-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bbd",
     9 => x"8c080b0b",
    10 => x"0bbd9008",
    11 => x"0b0b0bbd",
    12 => x"94080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"bd940c0b",
    16 => x"0b0bbd90",
    17 => x"0c0b0b0b",
    18 => x"bd8c0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb6d4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"bd8c7080",
    57 => x"c7c4278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"5188c204",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bbd9c0c",
    65 => x"9f0bbda0",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"bda008ff",
    69 => x"05bda00c",
    70 => x"bda00880",
    71 => x"25eb38bd",
    72 => x"9c08ff05",
    73 => x"bd9c0cbd",
    74 => x"9c088025",
    75 => x"d738800b",
    76 => x"bda00c80",
    77 => x"0bbd9c0c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bbd9c08",
    97 => x"258f3882",
    98 => x"bd2dbd9c",
    99 => x"08ff05bd",
   100 => x"9c0c82ff",
   101 => x"04bd9c08",
   102 => x"bda00853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"bd9c08a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134bda0",
   111 => x"088105bd",
   112 => x"a00cbda0",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bbda00c",
   116 => x"bd9c0881",
   117 => x"05bd9c0c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134bd",
   122 => x"a0088105",
   123 => x"bda00cbd",
   124 => x"a008a02e",
   125 => x"0981068e",
   126 => x"38800bbd",
   127 => x"a00cbd9c",
   128 => x"088105bd",
   129 => x"9c0c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bbda4",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bbda40c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872bd",
   169 => x"a4088407",
   170 => x"bda40c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb9b8",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"bda40852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"bd8c0c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c028405",
   216 => x"0d0402fc",
   217 => x"050dbde0",
   218 => x"0880c007",
   219 => x"ed0c0284",
   220 => x"050d0402",
   221 => x"fc050dbd",
   222 => x"e0088180",
   223 => x"07ed0c02",
   224 => x"84050d04",
   225 => x"880bec0c",
   226 => x"86b72d04",
   227 => x"900bec0c",
   228 => x"86b72d04",
   229 => x"02dc050d",
   230 => x"80598784",
   231 => x"2d810bec",
   232 => x"0c7a52bd",
   233 => x"a851adf5",
   234 => x"2dbd8c08",
   235 => x"792e80ee",
   236 => x"38bdac08",
   237 => x"70f80c79",
   238 => x"ff125659",
   239 => x"5573792e",
   240 => x"8b388118",
   241 => x"74812a55",
   242 => x"5873f738",
   243 => x"f7185881",
   244 => x"59807525",
   245 => x"80c83877",
   246 => x"52735184",
   247 => x"8b2dbdfc",
   248 => x"52bda851",
   249 => x"b0b42dbd",
   250 => x"8c08802e",
   251 => x"9a38bdfc",
   252 => x"5783fc56",
   253 => x"76708405",
   254 => x"5808e80c",
   255 => x"fc165675",
   256 => x"8025f138",
   257 => x"888e04bd",
   258 => x"8c085984",
   259 => x"8055bda8",
   260 => x"51b0862d",
   261 => x"fc801581",
   262 => x"15555587",
   263 => x"d104840b",
   264 => x"ec0c7880",
   265 => x"2e8d38b9",
   266 => x"bc5190fd",
   267 => x"2d8ef42d",
   268 => x"88b904ba",
   269 => x"9c5190fd",
   270 => x"2d78bd8c",
   271 => x"0c02a405",
   272 => x"0d0402ec",
   273 => x"050d840b",
   274 => x"ec0c8ec2",
   275 => x"2d8b912d",
   276 => x"81f82d83",
   277 => x"538ea72d",
   278 => x"815184f0",
   279 => x"2dff1353",
   280 => x"728025f1",
   281 => x"38840bec",
   282 => x"0cb7ec51",
   283 => x"85fe2da4",
   284 => x"ea2dbd8c",
   285 => x"08802e82",
   286 => x"8338810b",
   287 => x"ec0cb6e4",
   288 => x"52bda851",
   289 => x"adf52dbd",
   290 => x"8c08802e",
   291 => x"80c738bd",
   292 => x"fc52bda8",
   293 => x"51b0b42d",
   294 => x"bd8c0880",
   295 => x"2eb738bd",
   296 => x"fc0b80f5",
   297 => x"2dbbac0c",
   298 => x"bdfd0b80",
   299 => x"f52dbbb0",
   300 => x"0cbdfe0b",
   301 => x"80f52dbb",
   302 => x"b40cbdff",
   303 => x"0b80f52d",
   304 => x"bbb80cbe",
   305 => x"800b80f5",
   306 => x"2dbbbc0c",
   307 => x"be810b80",
   308 => x"f52dbbc0",
   309 => x"0cb6f452",
   310 => x"bda851ad",
   311 => x"f52dbd8c",
   312 => x"08802e80",
   313 => x"c738bdfc",
   314 => x"52bda851",
   315 => x"b0b42dbd",
   316 => x"8c08802e",
   317 => x"b738bdfc",
   318 => x"0b80f52d",
   319 => x"bb8c0cbd",
   320 => x"fd0b80f5",
   321 => x"2dbb900c",
   322 => x"bdfe0b80",
   323 => x"f52dbb94",
   324 => x"0cbdff0b",
   325 => x"80f52dbb",
   326 => x"980cbe80",
   327 => x"0b80f52d",
   328 => x"bb9c0cbe",
   329 => x"810b80f5",
   330 => x"2dbba00c",
   331 => x"879451b6",
   332 => x"ce2db9bc",
   333 => x"5190fd2d",
   334 => x"8ee12d8b",
   335 => x"9d2d918d",
   336 => x"2db9d00b",
   337 => x"80f52dbb",
   338 => x"88087081",
   339 => x"06555654",
   340 => x"72802e85",
   341 => x"38738107",
   342 => x"5474812a",
   343 => x"70810651",
   344 => x"5372802e",
   345 => x"85387382",
   346 => x"075473fc",
   347 => x"0c8653bd",
   348 => x"8c088338",
   349 => x"845372ec",
   350 => x"0c8abb04",
   351 => x"800bbd8c",
   352 => x"0c029405",
   353 => x"0d047198",
   354 => x"0c04ffb0",
   355 => x"08bd8c0c",
   356 => x"04810bff",
   357 => x"b00c0480",
   358 => x"0bffb00c",
   359 => x"0402f405",
   360 => x"0d8c9f04",
   361 => x"bd8c0881",
   362 => x"f02e0981",
   363 => x"06893881",
   364 => x"0bbb800c",
   365 => x"8c9f04bd",
   366 => x"8c0881e0",
   367 => x"2e098106",
   368 => x"8938810b",
   369 => x"bb840c8c",
   370 => x"9f04bd8c",
   371 => x"0852bb84",
   372 => x"08802e88",
   373 => x"38bd8c08",
   374 => x"81800552",
   375 => x"71842c72",
   376 => x"8f065353",
   377 => x"bb800880",
   378 => x"2e993872",
   379 => x"8429bac0",
   380 => x"05721381",
   381 => x"712b7009",
   382 => x"73080673",
   383 => x"0c515353",
   384 => x"8c950472",
   385 => x"8429bac0",
   386 => x"05721383",
   387 => x"712b7208",
   388 => x"07720c53",
   389 => x"53800bbb",
   390 => x"840c800b",
   391 => x"bb800cbd",
   392 => x"b4518da0",
   393 => x"2dbd8c08",
   394 => x"ff24fef8",
   395 => x"38800bbd",
   396 => x"8c0c028c",
   397 => x"050d0402",
   398 => x"f8050dba",
   399 => x"c0528f51",
   400 => x"80727084",
   401 => x"05540cff",
   402 => x"11517080",
   403 => x"25f23802",
   404 => x"88050d04",
   405 => x"02f0050d",
   406 => x"75518b97",
   407 => x"2d70822c",
   408 => x"fc06bac0",
   409 => x"1172109e",
   410 => x"06710870",
   411 => x"722a7083",
   412 => x"0682742b",
   413 => x"70097406",
   414 => x"760c5451",
   415 => x"56575351",
   416 => x"538b912d",
   417 => x"71bd8c0c",
   418 => x"0290050d",
   419 => x"0402fc05",
   420 => x"0d725180",
   421 => x"710c800b",
   422 => x"84120c02",
   423 => x"84050d04",
   424 => x"02f0050d",
   425 => x"75700884",
   426 => x"12085353",
   427 => x"53ff5471",
   428 => x"712ea838",
   429 => x"8b972d84",
   430 => x"13087084",
   431 => x"29148811",
   432 => x"70087081",
   433 => x"ff068418",
   434 => x"08811187",
   435 => x"06841a0c",
   436 => x"53515551",
   437 => x"51518b91",
   438 => x"2d715473",
   439 => x"bd8c0c02",
   440 => x"90050d04",
   441 => x"02f8050d",
   442 => x"8b972de0",
   443 => x"08708b2a",
   444 => x"70810651",
   445 => x"52527080",
   446 => x"2e9d38bd",
   447 => x"b4087084",
   448 => x"29bdbc05",
   449 => x"7381ff06",
   450 => x"710c5151",
   451 => x"bdb40881",
   452 => x"118706bd",
   453 => x"b40c5180",
   454 => x"0bbddc0c",
   455 => x"8b8a2d8b",
   456 => x"912d0288",
   457 => x"050d0402",
   458 => x"fc050d8b",
   459 => x"972d810b",
   460 => x"bddc0c8b",
   461 => x"912dbddc",
   462 => x"085170fa",
   463 => x"38028405",
   464 => x"0d0402fc",
   465 => x"050dbdb4",
   466 => x"518d8d2d",
   467 => x"8cb72d8d",
   468 => x"e4518b86",
   469 => x"2d028405",
   470 => x"0d04bde8",
   471 => x"08bd8c0c",
   472 => x"0402fc05",
   473 => x"0d810bbb",
   474 => x"cc0c8151",
   475 => x"84f02d02",
   476 => x"84050d04",
   477 => x"02fc050d",
   478 => x"8efe048b",
   479 => x"9d2d80f6",
   480 => x"518cd42d",
   481 => x"bd8c08f3",
   482 => x"3880da51",
   483 => x"8cd42dbd",
   484 => x"8c08e838",
   485 => x"bbbc0851",
   486 => x"8cd42dbd",
   487 => x"8c08dc38",
   488 => x"bd8c08bb",
   489 => x"cc0cbd8c",
   490 => x"085184f0",
   491 => x"2d028405",
   492 => x"0d0402ec",
   493 => x"050d7654",
   494 => x"8052870b",
   495 => x"881580f5",
   496 => x"2d565374",
   497 => x"72248338",
   498 => x"a0537251",
   499 => x"82f92d81",
   500 => x"128b1580",
   501 => x"f52d5452",
   502 => x"727225de",
   503 => x"38029405",
   504 => x"0d0402f0",
   505 => x"050dbde8",
   506 => x"085481f8",
   507 => x"2d800bbd",
   508 => x"ec0c7308",
   509 => x"802e8180",
   510 => x"38820bbd",
   511 => x"a00cbdec",
   512 => x"088f06bd",
   513 => x"9c0c7308",
   514 => x"5271832e",
   515 => x"96387183",
   516 => x"26893871",
   517 => x"812eaf38",
   518 => x"90e30471",
   519 => x"852e9f38",
   520 => x"90e30488",
   521 => x"1480f52d",
   522 => x"841508b8",
   523 => x"84535452",
   524 => x"85fe2d71",
   525 => x"84291370",
   526 => x"08525290",
   527 => x"e7047351",
   528 => x"8fb22d90",
   529 => x"e304bb88",
   530 => x"08881508",
   531 => x"2c708106",
   532 => x"51527180",
   533 => x"2e8738b8",
   534 => x"885190e0",
   535 => x"04b88c51",
   536 => x"85fe2d84",
   537 => x"14085185",
   538 => x"fe2dbdec",
   539 => x"088105bd",
   540 => x"ec0c8c14",
   541 => x"548ff204",
   542 => x"0290050d",
   543 => x"0471bde8",
   544 => x"0c8fe22d",
   545 => x"bdec08ff",
   546 => x"05bdf00c",
   547 => x"0402e805",
   548 => x"0dbde808",
   549 => x"bdf40857",
   550 => x"5580f651",
   551 => x"8cd42dbd",
   552 => x"8c08812a",
   553 => x"70810651",
   554 => x"5271802e",
   555 => x"9f3891b4",
   556 => x"048b9d2d",
   557 => x"80f6518c",
   558 => x"d42dbd8c",
   559 => x"08f338bb",
   560 => x"cc088132",
   561 => x"70bbcc0c",
   562 => x"5184f02d",
   563 => x"800bbde0",
   564 => x"0c800bbd",
   565 => x"e40c8c51",
   566 => x"8cd42dbd",
   567 => x"8c08812a",
   568 => x"70810651",
   569 => x"5271802e",
   570 => x"80e338bb",
   571 => x"8c08bbac",
   572 => x"08bb8c0c",
   573 => x"bbac0cbb",
   574 => x"9008bbb0",
   575 => x"08bb900c",
   576 => x"bbb00cbb",
   577 => x"9408bbb4",
   578 => x"08bb940c",
   579 => x"bbb40cbb",
   580 => x"9808bbb8",
   581 => x"08bb980c",
   582 => x"bbb80cbb",
   583 => x"9c08bbbc",
   584 => x"08bb9c0c",
   585 => x"bbbc0cbb",
   586 => x"a008bbc0",
   587 => x"08bba00c",
   588 => x"bbc00cbb",
   589 => x"a408bbc4",
   590 => x"08bba40c",
   591 => x"bbc40cbb",
   592 => x"a808bbc8",
   593 => x"08bba80c",
   594 => x"70bbc80c",
   595 => x"52bbcc08",
   596 => x"83bc38bb",
   597 => x"ac08518c",
   598 => x"d42dbd8c",
   599 => x"08802e89",
   600 => x"38bde008",
   601 => x"8107bde0",
   602 => x"0cbbb008",
   603 => x"518cd42d",
   604 => x"bd8c0880",
   605 => x"2e8938bd",
   606 => x"e0088207",
   607 => x"bde00cbb",
   608 => x"b408518c",
   609 => x"d42dbd8c",
   610 => x"08802e89",
   611 => x"38bde008",
   612 => x"8407bde0",
   613 => x"0cbbb808",
   614 => x"518cd42d",
   615 => x"bd8c0880",
   616 => x"2e8938bd",
   617 => x"e0088807",
   618 => x"bde00cbb",
   619 => x"bc08518c",
   620 => x"d42dbd8c",
   621 => x"08802e89",
   622 => x"38bde008",
   623 => x"9007bde0",
   624 => x"0cbbc008",
   625 => x"518cd42d",
   626 => x"bd8c0880",
   627 => x"2e8938bd",
   628 => x"e008a007",
   629 => x"bde00cbb",
   630 => x"c408518c",
   631 => x"d42dbd8c",
   632 => x"08802e8a",
   633 => x"38bde008",
   634 => x"80c007bd",
   635 => x"e00cbbc8",
   636 => x"08518cd4",
   637 => x"2dbd8c08",
   638 => x"802e8a38",
   639 => x"bde00881",
   640 => x"8007bde0",
   641 => x"0cbb8c08",
   642 => x"518cd42d",
   643 => x"bd8c0880",
   644 => x"2e8938bd",
   645 => x"e4088107",
   646 => x"bde40cbb",
   647 => x"9008518c",
   648 => x"d42dbd8c",
   649 => x"08802e89",
   650 => x"38bde408",
   651 => x"8207bde4",
   652 => x"0cbb9408",
   653 => x"518cd42d",
   654 => x"bd8c0880",
   655 => x"2e8938bd",
   656 => x"e4088407",
   657 => x"bde40cbb",
   658 => x"9808518c",
   659 => x"d42dbd8c",
   660 => x"08802e89",
   661 => x"38bde408",
   662 => x"8807bde4",
   663 => x"0cbb9c08",
   664 => x"518cd42d",
   665 => x"bd8c0880",
   666 => x"2e8938bd",
   667 => x"e4089007",
   668 => x"bde40cbb",
   669 => x"a008518c",
   670 => x"d42dbd8c",
   671 => x"08802e89",
   672 => x"38bde408",
   673 => x"a007bde4",
   674 => x"0cbba408",
   675 => x"518cd42d",
   676 => x"bd8c0880",
   677 => x"2e8a38bd",
   678 => x"e40880c0",
   679 => x"07bde40c",
   680 => x"bba80851",
   681 => x"8cd42dbd",
   682 => x"8c08802e",
   683 => x"8a38bde4",
   684 => x"08818007",
   685 => x"bde40cbd",
   686 => x"e008ed0c",
   687 => x"bde408ee",
   688 => x"0c94518c",
   689 => x"d42dbd8c",
   690 => x"088e3881",
   691 => x"94518cd4",
   692 => x"2dbd8c08",
   693 => x"802ea838",
   694 => x"91518cd4",
   695 => x"2dbd8c08",
   696 => x"8e388191",
   697 => x"518cd42d",
   698 => x"bd8c0880",
   699 => x"2e913880",
   700 => x"e6518cd4",
   701 => x"2dbd8c08",
   702 => x"802e8438",
   703 => x"878c2d81",
   704 => x"fd518cd4",
   705 => x"2d81fa51",
   706 => x"8cd42d9c",
   707 => x"e1049451",
   708 => x"8cd42dbd",
   709 => x"8c088e38",
   710 => x"8194518c",
   711 => x"d42dbd8c",
   712 => x"08802ea8",
   713 => x"3891518c",
   714 => x"d42dbd8c",
   715 => x"088e3881",
   716 => x"91518cd4",
   717 => x"2dbd8c08",
   718 => x"802e9138",
   719 => x"80e6518c",
   720 => x"d42dbd8c",
   721 => x"08802e84",
   722 => x"38878c2d",
   723 => x"81f5518c",
   724 => x"d42dbd8c",
   725 => x"08812a70",
   726 => x"81065152",
   727 => x"719738bb",
   728 => x"ac08518c",
   729 => x"d42dbd8c",
   730 => x"08812a70",
   731 => x"81065152",
   732 => x"71802eaf",
   733 => x"38bdf008",
   734 => x"5271802e",
   735 => x"8938ff12",
   736 => x"bdf00c97",
   737 => x"a304bdec",
   738 => x"0810bdec",
   739 => x"08057084",
   740 => x"29165152",
   741 => x"88120880",
   742 => x"2e8938ff",
   743 => x"51881208",
   744 => x"52712d81",
   745 => x"f2518cd4",
   746 => x"2dbd8c08",
   747 => x"812a7081",
   748 => x"06515271",
   749 => x"9738bbb0",
   750 => x"08518cd4",
   751 => x"2dbd8c08",
   752 => x"812a7081",
   753 => x"06515271",
   754 => x"802eb138",
   755 => x"bdec08ff",
   756 => x"11bdf008",
   757 => x"56535373",
   758 => x"72258938",
   759 => x"8114bdf0",
   760 => x"0c97fc04",
   761 => x"72101370",
   762 => x"84291651",
   763 => x"52881208",
   764 => x"802e8938",
   765 => x"fe518812",
   766 => x"0852712d",
   767 => x"81fd518c",
   768 => x"d42dbd8c",
   769 => x"08812a70",
   770 => x"81065152",
   771 => x"719738bb",
   772 => x"b408518c",
   773 => x"d42dbd8c",
   774 => x"08812a70",
   775 => x"81065152",
   776 => x"71802ead",
   777 => x"38bdf008",
   778 => x"802e8938",
   779 => x"800bbdf0",
   780 => x"0c98d104",
   781 => x"bdec0810",
   782 => x"bdec0805",
   783 => x"70842916",
   784 => x"51528812",
   785 => x"08802e89",
   786 => x"38fd5188",
   787 => x"12085271",
   788 => x"2d81fa51",
   789 => x"8cd42dbd",
   790 => x"8c08812a",
   791 => x"70810651",
   792 => x"52719738",
   793 => x"bbb80851",
   794 => x"8cd42dbd",
   795 => x"8c08812a",
   796 => x"70810651",
   797 => x"5271802e",
   798 => x"ae38bdec",
   799 => x"08ff1154",
   800 => x"52bdf008",
   801 => x"73258838",
   802 => x"72bdf00c",
   803 => x"99a70471",
   804 => x"10127084",
   805 => x"29165152",
   806 => x"88120880",
   807 => x"2e8938fc",
   808 => x"51881208",
   809 => x"52712dbd",
   810 => x"f0087053",
   811 => x"5473802e",
   812 => x"8a388c15",
   813 => x"ff155555",
   814 => x"99ad0482",
   815 => x"0bbda00c",
   816 => x"718f06bd",
   817 => x"9c0c81eb",
   818 => x"518cd42d",
   819 => x"bd8c0881",
   820 => x"2a708106",
   821 => x"51527180",
   822 => x"2ead3874",
   823 => x"08852e09",
   824 => x"8106a438",
   825 => x"881580f5",
   826 => x"2dff0552",
   827 => x"71881681",
   828 => x"b72d7198",
   829 => x"2b527180",
   830 => x"25883880",
   831 => x"0b881681",
   832 => x"b72d7451",
   833 => x"8fb22d81",
   834 => x"f4518cd4",
   835 => x"2dbd8c08",
   836 => x"812a7081",
   837 => x"06515271",
   838 => x"802eb338",
   839 => x"7408852e",
   840 => x"098106aa",
   841 => x"38881580",
   842 => x"f52d8105",
   843 => x"52718816",
   844 => x"81b72d71",
   845 => x"81ff068b",
   846 => x"1680f52d",
   847 => x"54527272",
   848 => x"27873872",
   849 => x"881681b7",
   850 => x"2d74518f",
   851 => x"b22d80da",
   852 => x"518cd42d",
   853 => x"bd8c0881",
   854 => x"2a708106",
   855 => x"51527198",
   856 => x"38bbbc08",
   857 => x"518cd42d",
   858 => x"bd8c0881",
   859 => x"2a708106",
   860 => x"51527180",
   861 => x"2e81a638",
   862 => x"bde808bd",
   863 => x"f0085553",
   864 => x"73802e8a",
   865 => x"388c13ff",
   866 => x"1555539b",
   867 => x"80047208",
   868 => x"5271822e",
   869 => x"a6387182",
   870 => x"26893871",
   871 => x"812ea938",
   872 => x"9c9d0471",
   873 => x"832eb138",
   874 => x"71842e09",
   875 => x"810680ed",
   876 => x"38881308",
   877 => x"5190fd2d",
   878 => x"9c9d04bd",
   879 => x"f0085188",
   880 => x"13085271",
   881 => x"2d9c9d04",
   882 => x"810b8814",
   883 => x"082bbb88",
   884 => x"0832bb88",
   885 => x"0c9bf304",
   886 => x"881380f5",
   887 => x"2d81058b",
   888 => x"1480f52d",
   889 => x"53547174",
   890 => x"24833880",
   891 => x"54738814",
   892 => x"81b72d8f",
   893 => x"e22d9c9d",
   894 => x"04750880",
   895 => x"2ea23875",
   896 => x"08518cd4",
   897 => x"2dbd8c08",
   898 => x"81065271",
   899 => x"802e8b38",
   900 => x"bdf00851",
   901 => x"84160852",
   902 => x"712d8816",
   903 => x"5675da38",
   904 => x"8054800b",
   905 => x"bda00c73",
   906 => x"8f06bd9c",
   907 => x"0ca05273",
   908 => x"bdf0082e",
   909 => x"09810698",
   910 => x"38bdec08",
   911 => x"ff057432",
   912 => x"70098105",
   913 => x"7072079f",
   914 => x"2a917131",
   915 => x"51515353",
   916 => x"715182f9",
   917 => x"2d811454",
   918 => x"8e7425c6",
   919 => x"38bbcc08",
   920 => x"5271bd8c",
   921 => x"0c029805",
   922 => x"0d0402f4",
   923 => x"050dd452",
   924 => x"81ff720c",
   925 => x"71085381",
   926 => x"ff720c72",
   927 => x"882b83fe",
   928 => x"80067208",
   929 => x"7081ff06",
   930 => x"51525381",
   931 => x"ff720c72",
   932 => x"7107882b",
   933 => x"72087081",
   934 => x"ff065152",
   935 => x"5381ff72",
   936 => x"0c727107",
   937 => x"882b7208",
   938 => x"7081ff06",
   939 => x"7207bd8c",
   940 => x"0c525302",
   941 => x"8c050d04",
   942 => x"02f4050d",
   943 => x"74767181",
   944 => x"ff06d40c",
   945 => x"5353bdf8",
   946 => x"08853871",
   947 => x"892b5271",
   948 => x"982ad40c",
   949 => x"71902a70",
   950 => x"81ff06d4",
   951 => x"0c517188",
   952 => x"2a7081ff",
   953 => x"06d40c51",
   954 => x"7181ff06",
   955 => x"d40c7290",
   956 => x"2a7081ff",
   957 => x"06d40c51",
   958 => x"d4087081",
   959 => x"ff065151",
   960 => x"82b8bf52",
   961 => x"7081ff2e",
   962 => x"09810694",
   963 => x"3881ff0b",
   964 => x"d40cd408",
   965 => x"7081ff06",
   966 => x"ff145451",
   967 => x"5171e538",
   968 => x"70bd8c0c",
   969 => x"028c050d",
   970 => x"0402fc05",
   971 => x"0d81c751",
   972 => x"81ff0bd4",
   973 => x"0cff1151",
   974 => x"708025f4",
   975 => x"38028405",
   976 => x"0d0402f4",
   977 => x"050d81ff",
   978 => x"0bd40c93",
   979 => x"53805287",
   980 => x"fc80c151",
   981 => x"9db82dbd",
   982 => x"8c088b38",
   983 => x"81ff0bd4",
   984 => x"0c81539e",
   985 => x"ef049ea9",
   986 => x"2dff1353",
   987 => x"72df3872",
   988 => x"bd8c0c02",
   989 => x"8c050d04",
   990 => x"02ec050d",
   991 => x"810bbdf8",
   992 => x"0c8454d0",
   993 => x"08708f2a",
   994 => x"70810651",
   995 => x"515372f3",
   996 => x"3872d00c",
   997 => x"9ea92db8",
   998 => x"905185fe",
   999 => x"2dd00870",
  1000 => x"8f2a7081",
  1001 => x"06515153",
  1002 => x"72f33881",
  1003 => x"0bd00cb1",
  1004 => x"53805284",
  1005 => x"d480c051",
  1006 => x"9db82dbd",
  1007 => x"8c08812e",
  1008 => x"93387282",
  1009 => x"2ebd38ff",
  1010 => x"135372e5",
  1011 => x"38ff1454",
  1012 => x"73ffb038",
  1013 => x"9ea92d83",
  1014 => x"aa52849c",
  1015 => x"80c8519d",
  1016 => x"b82dbd8c",
  1017 => x"08812e09",
  1018 => x"81069238",
  1019 => x"9cea2dbd",
  1020 => x"8c0883ff",
  1021 => x"ff065372",
  1022 => x"83aa2e9d",
  1023 => x"389ec22d",
  1024 => x"a09404b8",
  1025 => x"9c5185fe",
  1026 => x"2d8053a1",
  1027 => x"e204b8b4",
  1028 => x"5185fe2d",
  1029 => x"8054a1b4",
  1030 => x"0481ff0b",
  1031 => x"d40cb154",
  1032 => x"9ea92d8f",
  1033 => x"cf538052",
  1034 => x"87fc80f7",
  1035 => x"519db82d",
  1036 => x"bd8c0855",
  1037 => x"bd8c0881",
  1038 => x"2e098106",
  1039 => x"9b3881ff",
  1040 => x"0bd40c82",
  1041 => x"0a52849c",
  1042 => x"80e9519d",
  1043 => x"b82dbd8c",
  1044 => x"08802e8d",
  1045 => x"389ea92d",
  1046 => x"ff135372",
  1047 => x"c938a1a7",
  1048 => x"0481ff0b",
  1049 => x"d40cbd8c",
  1050 => x"085287fc",
  1051 => x"80fa519d",
  1052 => x"b82dbd8c",
  1053 => x"08b13881",
  1054 => x"ff0bd40c",
  1055 => x"d4085381",
  1056 => x"ff0bd40c",
  1057 => x"81ff0bd4",
  1058 => x"0c81ff0b",
  1059 => x"d40c81ff",
  1060 => x"0bd40c72",
  1061 => x"862a7081",
  1062 => x"06765651",
  1063 => x"53729538",
  1064 => x"bd8c0854",
  1065 => x"a1b40473",
  1066 => x"822efee2",
  1067 => x"38ff1454",
  1068 => x"73feed38",
  1069 => x"73bdf80c",
  1070 => x"738b3881",
  1071 => x"5287fc80",
  1072 => x"d0519db8",
  1073 => x"2d81ff0b",
  1074 => x"d40cd008",
  1075 => x"708f2a70",
  1076 => x"81065151",
  1077 => x"5372f338",
  1078 => x"72d00c81",
  1079 => x"ff0bd40c",
  1080 => x"815372bd",
  1081 => x"8c0c0294",
  1082 => x"050d0402",
  1083 => x"e8050d78",
  1084 => x"55805681",
  1085 => x"ff0bd40c",
  1086 => x"d008708f",
  1087 => x"2a708106",
  1088 => x"51515372",
  1089 => x"f3388281",
  1090 => x"0bd00c81",
  1091 => x"ff0bd40c",
  1092 => x"775287fc",
  1093 => x"80d1519d",
  1094 => x"b82d80db",
  1095 => x"c6df54bd",
  1096 => x"8c08802e",
  1097 => x"8a38b8d4",
  1098 => x"5185fe2d",
  1099 => x"a3820481",
  1100 => x"ff0bd40c",
  1101 => x"d4087081",
  1102 => x"ff065153",
  1103 => x"7281fe2e",
  1104 => x"0981069d",
  1105 => x"3880ff53",
  1106 => x"9cea2dbd",
  1107 => x"8c087570",
  1108 => x"8405570c",
  1109 => x"ff135372",
  1110 => x"8025ed38",
  1111 => x"8156a2e7",
  1112 => x"04ff1454",
  1113 => x"73c93881",
  1114 => x"ff0bd40c",
  1115 => x"81ff0bd4",
  1116 => x"0cd00870",
  1117 => x"8f2a7081",
  1118 => x"06515153",
  1119 => x"72f33872",
  1120 => x"d00c75bd",
  1121 => x"8c0c0298",
  1122 => x"050d0402",
  1123 => x"e8050d77",
  1124 => x"797b5855",
  1125 => x"55805372",
  1126 => x"7625a338",
  1127 => x"74708105",
  1128 => x"5680f52d",
  1129 => x"74708105",
  1130 => x"5680f52d",
  1131 => x"52527171",
  1132 => x"2e863881",
  1133 => x"51a3c004",
  1134 => x"811353a3",
  1135 => x"97048051",
  1136 => x"70bd8c0c",
  1137 => x"0298050d",
  1138 => x"0402ec05",
  1139 => x"0d765574",
  1140 => x"802ebe38",
  1141 => x"9a1580e0",
  1142 => x"2d51b18d",
  1143 => x"2dbd8c08",
  1144 => x"bd8c0880",
  1145 => x"c4ac0cbd",
  1146 => x"8c085454",
  1147 => x"80c48808",
  1148 => x"802e9938",
  1149 => x"941580e0",
  1150 => x"2d51b18d",
  1151 => x"2dbd8c08",
  1152 => x"902b83ff",
  1153 => x"f00a0670",
  1154 => x"75075153",
  1155 => x"7280c4ac",
  1156 => x"0c80c4ac",
  1157 => x"08537280",
  1158 => x"2e9d3880",
  1159 => x"c48008fe",
  1160 => x"14712980",
  1161 => x"c4940805",
  1162 => x"80c4b00c",
  1163 => x"70842b80",
  1164 => x"c48c0c54",
  1165 => x"a4e50480",
  1166 => x"c4980880",
  1167 => x"c4ac0c80",
  1168 => x"c49c0880",
  1169 => x"c4b00c80",
  1170 => x"c4880880",
  1171 => x"2e8b3880",
  1172 => x"c4800884",
  1173 => x"2b53a4e0",
  1174 => x"0480c4a0",
  1175 => x"08842b53",
  1176 => x"7280c48c",
  1177 => x"0c029405",
  1178 => x"0d0402d8",
  1179 => x"050d800b",
  1180 => x"80c4880c",
  1181 => x"84549ef8",
  1182 => x"2dbd8c08",
  1183 => x"802e9538",
  1184 => x"bdfc5280",
  1185 => x"51a1eb2d",
  1186 => x"bd8c0880",
  1187 => x"2e8638fe",
  1188 => x"54a59c04",
  1189 => x"ff145473",
  1190 => x"8024db38",
  1191 => x"738c38b8",
  1192 => x"e45185fe",
  1193 => x"2d7355aa",
  1194 => x"c6048056",
  1195 => x"810b80c4",
  1196 => x"b40c8853",
  1197 => x"b8f852be",
  1198 => x"b251a38b",
  1199 => x"2dbd8c08",
  1200 => x"762e0981",
  1201 => x"068838bd",
  1202 => x"8c0880c4",
  1203 => x"b40c8853",
  1204 => x"b98452be",
  1205 => x"ce51a38b",
  1206 => x"2dbd8c08",
  1207 => x"8838bd8c",
  1208 => x"0880c4b4",
  1209 => x"0c80c4b4",
  1210 => x"08802e80",
  1211 => x"fc3880c1",
  1212 => x"c20b80f5",
  1213 => x"2d80c1c3",
  1214 => x"0b80f52d",
  1215 => x"71982b71",
  1216 => x"902b0780",
  1217 => x"c1c40b80",
  1218 => x"f52d7088",
  1219 => x"2b720780",
  1220 => x"c1c50b80",
  1221 => x"f52d7107",
  1222 => x"80c1fa0b",
  1223 => x"80f52d80",
  1224 => x"c1fb0b80",
  1225 => x"f52d7188",
  1226 => x"2b07535f",
  1227 => x"54525a56",
  1228 => x"57557381",
  1229 => x"abaa2e09",
  1230 => x"81068d38",
  1231 => x"7551b0dd",
  1232 => x"2dbd8c08",
  1233 => x"56a6d504",
  1234 => x"7382d4d5",
  1235 => x"2e8738b9",
  1236 => x"9051a797",
  1237 => x"04bdfc52",
  1238 => x"7551a1eb",
  1239 => x"2dbd8c08",
  1240 => x"55bd8c08",
  1241 => x"802e83de",
  1242 => x"388853b9",
  1243 => x"8452bece",
  1244 => x"51a38b2d",
  1245 => x"bd8c088a",
  1246 => x"38810b80",
  1247 => x"c4880ca7",
  1248 => x"9d048853",
  1249 => x"b8f852be",
  1250 => x"b251a38b",
  1251 => x"2dbd8c08",
  1252 => x"802e8a38",
  1253 => x"b9a45185",
  1254 => x"fe2da7f9",
  1255 => x"0480c1fa",
  1256 => x"0b80f52d",
  1257 => x"547380d5",
  1258 => x"2e098106",
  1259 => x"80cb3880",
  1260 => x"c1fb0b80",
  1261 => x"f52d5473",
  1262 => x"81aa2e09",
  1263 => x"8106ba38",
  1264 => x"800bbdfc",
  1265 => x"0b80f52d",
  1266 => x"56547481",
  1267 => x"e92e8338",
  1268 => x"81547481",
  1269 => x"eb2e8c38",
  1270 => x"80557375",
  1271 => x"2e098106",
  1272 => x"82e438be",
  1273 => x"870b80f5",
  1274 => x"2d55748d",
  1275 => x"38be880b",
  1276 => x"80f52d54",
  1277 => x"73822e86",
  1278 => x"388055aa",
  1279 => x"c604be89",
  1280 => x"0b80f52d",
  1281 => x"7080c480",
  1282 => x"0cff0580",
  1283 => x"c4840cbe",
  1284 => x"8a0b80f5",
  1285 => x"2dbe8b0b",
  1286 => x"80f52d58",
  1287 => x"76057782",
  1288 => x"80290570",
  1289 => x"80c4900c",
  1290 => x"be8c0b80",
  1291 => x"f52d7080",
  1292 => x"c4a40c80",
  1293 => x"c4880859",
  1294 => x"57587680",
  1295 => x"2e81ac38",
  1296 => x"8853b984",
  1297 => x"52bece51",
  1298 => x"a38b2dbd",
  1299 => x"8c0881f6",
  1300 => x"3880c480",
  1301 => x"0870842b",
  1302 => x"80c48c0c",
  1303 => x"7080c4a0",
  1304 => x"0cbea10b",
  1305 => x"80f52dbe",
  1306 => x"a00b80f5",
  1307 => x"2d718280",
  1308 => x"2905bea2",
  1309 => x"0b80f52d",
  1310 => x"70848080",
  1311 => x"2912bea3",
  1312 => x"0b80f52d",
  1313 => x"7081800a",
  1314 => x"29127080",
  1315 => x"c4a80c80",
  1316 => x"c4a40871",
  1317 => x"2980c490",
  1318 => x"08057080",
  1319 => x"c4940cbe",
  1320 => x"a90b80f5",
  1321 => x"2dbea80b",
  1322 => x"80f52d71",
  1323 => x"82802905",
  1324 => x"beaa0b80",
  1325 => x"f52d7084",
  1326 => x"80802912",
  1327 => x"beab0b80",
  1328 => x"f52d7098",
  1329 => x"2b81f00a",
  1330 => x"06720570",
  1331 => x"80c4980c",
  1332 => x"fe117e29",
  1333 => x"770580c4",
  1334 => x"9c0c5259",
  1335 => x"5243545e",
  1336 => x"51525952",
  1337 => x"5d575957",
  1338 => x"aabf04be",
  1339 => x"8e0b80f5",
  1340 => x"2dbe8d0b",
  1341 => x"80f52d71",
  1342 => x"82802905",
  1343 => x"7080c48c",
  1344 => x"0c70a029",
  1345 => x"83ff0570",
  1346 => x"892a7080",
  1347 => x"c4a00cbe",
  1348 => x"930b80f5",
  1349 => x"2dbe920b",
  1350 => x"80f52d71",
  1351 => x"82802905",
  1352 => x"7080c4a8",
  1353 => x"0c7b7129",
  1354 => x"1e7080c4",
  1355 => x"9c0c7d80",
  1356 => x"c4980c73",
  1357 => x"0580c494",
  1358 => x"0c555e51",
  1359 => x"51555580",
  1360 => x"51a3c92d",
  1361 => x"815574bd",
  1362 => x"8c0c02a8",
  1363 => x"050d0402",
  1364 => x"ec050d76",
  1365 => x"70872c71",
  1366 => x"80ff0655",
  1367 => x"565480c4",
  1368 => x"88088a38",
  1369 => x"73882c74",
  1370 => x"81ff0654",
  1371 => x"55bdfc52",
  1372 => x"80c49008",
  1373 => x"1551a1eb",
  1374 => x"2dbd8c08",
  1375 => x"54bd8c08",
  1376 => x"802eb438",
  1377 => x"80c48808",
  1378 => x"802e9838",
  1379 => x"728429bd",
  1380 => x"fc057008",
  1381 => x"5253b0dd",
  1382 => x"2dbd8c08",
  1383 => x"f00a0653",
  1384 => x"abb50472",
  1385 => x"10bdfc05",
  1386 => x"7080e02d",
  1387 => x"5253b18d",
  1388 => x"2dbd8c08",
  1389 => x"53725473",
  1390 => x"bd8c0c02",
  1391 => x"94050d04",
  1392 => x"02e0050d",
  1393 => x"7970842c",
  1394 => x"80c4b008",
  1395 => x"05718f06",
  1396 => x"52555372",
  1397 => x"8938bdfc",
  1398 => x"527351a1",
  1399 => x"eb2d72a0",
  1400 => x"29bdfc05",
  1401 => x"54807480",
  1402 => x"f52d5653",
  1403 => x"74732e83",
  1404 => x"38815374",
  1405 => x"81e52e81",
  1406 => x"f1388170",
  1407 => x"74065458",
  1408 => x"72802e81",
  1409 => x"e5388b14",
  1410 => x"80f52d70",
  1411 => x"832a7906",
  1412 => x"58567699",
  1413 => x"38bbd008",
  1414 => x"53728938",
  1415 => x"7280c1fc",
  1416 => x"0b81b72d",
  1417 => x"76bbd00c",
  1418 => x"7353adec",
  1419 => x"04758f2e",
  1420 => x"09810681",
  1421 => x"b538749f",
  1422 => x"068d2980",
  1423 => x"c1ef1151",
  1424 => x"53811480",
  1425 => x"f52d7370",
  1426 => x"81055581",
  1427 => x"b72d8314",
  1428 => x"80f52d73",
  1429 => x"70810555",
  1430 => x"81b72d85",
  1431 => x"1480f52d",
  1432 => x"73708105",
  1433 => x"5581b72d",
  1434 => x"871480f5",
  1435 => x"2d737081",
  1436 => x"055581b7",
  1437 => x"2d891480",
  1438 => x"f52d7370",
  1439 => x"81055581",
  1440 => x"b72d8e14",
  1441 => x"80f52d73",
  1442 => x"70810555",
  1443 => x"81b72d90",
  1444 => x"1480f52d",
  1445 => x"73708105",
  1446 => x"5581b72d",
  1447 => x"921480f5",
  1448 => x"2d737081",
  1449 => x"055581b7",
  1450 => x"2d941480",
  1451 => x"f52d7370",
  1452 => x"81055581",
  1453 => x"b72d9614",
  1454 => x"80f52d73",
  1455 => x"70810555",
  1456 => x"81b72d98",
  1457 => x"1480f52d",
  1458 => x"73708105",
  1459 => x"5581b72d",
  1460 => x"9c1480f5",
  1461 => x"2d737081",
  1462 => x"055581b7",
  1463 => x"2d9e1480",
  1464 => x"f52d7381",
  1465 => x"b72d77bb",
  1466 => x"d00c8053",
  1467 => x"72bd8c0c",
  1468 => x"02a0050d",
  1469 => x"0402cc05",
  1470 => x"0d7e605e",
  1471 => x"5a800b80",
  1472 => x"c4ac0880",
  1473 => x"c4b00859",
  1474 => x"5c568058",
  1475 => x"80c48c08",
  1476 => x"782e81b0",
  1477 => x"38778f06",
  1478 => x"a0175754",
  1479 => x"738f38bd",
  1480 => x"fc527651",
  1481 => x"811757a1",
  1482 => x"eb2dbdfc",
  1483 => x"56807680",
  1484 => x"f52d5654",
  1485 => x"74742e83",
  1486 => x"38815474",
  1487 => x"81e52e80",
  1488 => x"f7388170",
  1489 => x"7506555c",
  1490 => x"73802e80",
  1491 => x"eb388b16",
  1492 => x"80f52d98",
  1493 => x"06597880",
  1494 => x"df388b53",
  1495 => x"7c527551",
  1496 => x"a38b2dbd",
  1497 => x"8c0880d0",
  1498 => x"389c1608",
  1499 => x"51b0dd2d",
  1500 => x"bd8c0884",
  1501 => x"1b0c9a16",
  1502 => x"80e02d51",
  1503 => x"b18d2dbd",
  1504 => x"8c08bd8c",
  1505 => x"08881c0c",
  1506 => x"bd8c0855",
  1507 => x"5580c488",
  1508 => x"08802e98",
  1509 => x"38941680",
  1510 => x"e02d51b1",
  1511 => x"8d2dbd8c",
  1512 => x"08902b83",
  1513 => x"fff00a06",
  1514 => x"70165154",
  1515 => x"73881b0c",
  1516 => x"787a0c7b",
  1517 => x"54affd04",
  1518 => x"81185880",
  1519 => x"c48c0878",
  1520 => x"26fed238",
  1521 => x"80c48808",
  1522 => x"802eb038",
  1523 => x"7a51aacf",
  1524 => x"2dbd8c08",
  1525 => x"bd8c0880",
  1526 => x"fffffff8",
  1527 => x"06555b73",
  1528 => x"80ffffff",
  1529 => x"f82e9438",
  1530 => x"bd8c08fe",
  1531 => x"0580c480",
  1532 => x"082980c4",
  1533 => x"94080557",
  1534 => x"ae8a0480",
  1535 => x"5473bd8c",
  1536 => x"0c02b405",
  1537 => x"0d0402f4",
  1538 => x"050d7470",
  1539 => x"08810571",
  1540 => x"0c700880",
  1541 => x"c4840806",
  1542 => x"5353718e",
  1543 => x"38881308",
  1544 => x"51aacf2d",
  1545 => x"bd8c0888",
  1546 => x"140c810b",
  1547 => x"bd8c0c02",
  1548 => x"8c050d04",
  1549 => x"02f0050d",
  1550 => x"75881108",
  1551 => x"fe0580c4",
  1552 => x"80082980",
  1553 => x"c4940811",
  1554 => x"720880c4",
  1555 => x"84080605",
  1556 => x"79555354",
  1557 => x"54a1eb2d",
  1558 => x"0290050d",
  1559 => x"0402f405",
  1560 => x"0d747088",
  1561 => x"2a83fe80",
  1562 => x"06707298",
  1563 => x"2a077288",
  1564 => x"2b87fc80",
  1565 => x"80067398",
  1566 => x"2b81f00a",
  1567 => x"06717307",
  1568 => x"07bd8c0c",
  1569 => x"56515351",
  1570 => x"028c050d",
  1571 => x"0402f805",
  1572 => x"0d028e05",
  1573 => x"80f52d74",
  1574 => x"882b0770",
  1575 => x"83ffff06",
  1576 => x"bd8c0c51",
  1577 => x"0288050d",
  1578 => x"0402f405",
  1579 => x"0d747678",
  1580 => x"53545280",
  1581 => x"71259738",
  1582 => x"72708105",
  1583 => x"5480f52d",
  1584 => x"72708105",
  1585 => x"5481b72d",
  1586 => x"ff115170",
  1587 => x"eb388072",
  1588 => x"81b72d02",
  1589 => x"8c050d04",
  1590 => x"02e8050d",
  1591 => x"77568070",
  1592 => x"56547376",
  1593 => x"24b33880",
  1594 => x"c48c0874",
  1595 => x"2eab3873",
  1596 => x"51abc02d",
  1597 => x"bd8c08bd",
  1598 => x"8c080981",
  1599 => x"0570bd8c",
  1600 => x"08079f2a",
  1601 => x"77058117",
  1602 => x"57575353",
  1603 => x"74762489",
  1604 => x"3880c48c",
  1605 => x"087426d7",
  1606 => x"3872bd8c",
  1607 => x"0c029805",
  1608 => x"0d0402f0",
  1609 => x"050dbd88",
  1610 => x"081651b1",
  1611 => x"d82dbd8c",
  1612 => x"08802e9e",
  1613 => x"388b53bd",
  1614 => x"8c085280",
  1615 => x"c1fc51b1",
  1616 => x"a92d80c4",
  1617 => x"b8085473",
  1618 => x"802e8738",
  1619 => x"80c1fc51",
  1620 => x"732d0290",
  1621 => x"050d0402",
  1622 => x"dc050d80",
  1623 => x"705a5574",
  1624 => x"bd880825",
  1625 => x"b13880c4",
  1626 => x"8c08752e",
  1627 => x"a9387851",
  1628 => x"abc02dbd",
  1629 => x"8c080981",
  1630 => x"0570bd8c",
  1631 => x"08079f2a",
  1632 => x"7605811b",
  1633 => x"5b565474",
  1634 => x"bd880825",
  1635 => x"893880c4",
  1636 => x"8c087926",
  1637 => x"d9388055",
  1638 => x"7880c48c",
  1639 => x"082781d4",
  1640 => x"387851ab",
  1641 => x"c02dbd8c",
  1642 => x"08802e81",
  1643 => x"a838bd8c",
  1644 => x"088b0580",
  1645 => x"f52d7084",
  1646 => x"2a708106",
  1647 => x"77107884",
  1648 => x"2b80c1fc",
  1649 => x"0b80f52d",
  1650 => x"5c5c5351",
  1651 => x"55567380",
  1652 => x"2e80c938",
  1653 => x"7416822b",
  1654 => x"b5980bbb",
  1655 => x"dc120c54",
  1656 => x"77753110",
  1657 => x"80c4bc11",
  1658 => x"55569074",
  1659 => x"70810556",
  1660 => x"81b72da0",
  1661 => x"7481b72d",
  1662 => x"7681ff06",
  1663 => x"81165854",
  1664 => x"73802e8a",
  1665 => x"389c5380",
  1666 => x"c1fc52b4",
  1667 => x"94048b53",
  1668 => x"bd8c0852",
  1669 => x"80c4be16",
  1670 => x"51b4cd04",
  1671 => x"7416822b",
  1672 => x"b2a20bbb",
  1673 => x"dc120c54",
  1674 => x"7681ff06",
  1675 => x"81165854",
  1676 => x"73802e8a",
  1677 => x"389c5380",
  1678 => x"c1fc52b4",
  1679 => x"c4048b53",
  1680 => x"bd8c0852",
  1681 => x"77753110",
  1682 => x"80c4bc05",
  1683 => x"517655b1",
  1684 => x"a92db4e9",
  1685 => x"04749029",
  1686 => x"75317010",
  1687 => x"80c4bc05",
  1688 => x"5154bd8c",
  1689 => x"087481b7",
  1690 => x"2d811959",
  1691 => x"748b24a3",
  1692 => x"38b39804",
  1693 => x"74902975",
  1694 => x"31701080",
  1695 => x"c4bc058c",
  1696 => x"77315751",
  1697 => x"54807481",
  1698 => x"b72d9e14",
  1699 => x"ff165654",
  1700 => x"74f33802",
  1701 => x"a4050d04",
  1702 => x"02fc050d",
  1703 => x"bd880813",
  1704 => x"51b1d82d",
  1705 => x"bd8c0880",
  1706 => x"2e8838bd",
  1707 => x"8c0851a3",
  1708 => x"c92d800b",
  1709 => x"bd880cb2",
  1710 => x"d72d8fe2",
  1711 => x"2d028405",
  1712 => x"0d0402fc",
  1713 => x"050d7251",
  1714 => x"70fd2ead",
  1715 => x"3870fd24",
  1716 => x"8a3870fc",
  1717 => x"2e80c438",
  1718 => x"b6a30470",
  1719 => x"fe2eb138",
  1720 => x"70ff2e09",
  1721 => x"8106bc38",
  1722 => x"bd880851",
  1723 => x"70802eb3",
  1724 => x"38ff11bd",
  1725 => x"880cb6a3",
  1726 => x"04bd8808",
  1727 => x"f00570bd",
  1728 => x"880c5170",
  1729 => x"80259c38",
  1730 => x"800bbd88",
  1731 => x"0cb6a304",
  1732 => x"bd880881",
  1733 => x"05bd880c",
  1734 => x"b6a304bd",
  1735 => x"88089005",
  1736 => x"bd880cb2",
  1737 => x"d72d8fe2",
  1738 => x"2d028405",
  1739 => x"0d0402fc",
  1740 => x"050d800b",
  1741 => x"bd880cb2",
  1742 => x"d72d8eda",
  1743 => x"2dbd8c08",
  1744 => x"bcf80cbb",
  1745 => x"d45190fd",
  1746 => x"2d028405",
  1747 => x"0d047180",
  1748 => x"c4b80c04",
  1749 => x"00ffffff",
  1750 => x"ff00ffff",
  1751 => x"ffff00ff",
  1752 => x"ffffff00",
  1753 => x"4b455953",
  1754 => x"50312020",
  1755 => x"20202000",
  1756 => x"00000000",
  1757 => x"4b455953",
  1758 => x"50322020",
  1759 => x"20202000",
  1760 => x"00000000",
  1761 => x"52657365",
  1762 => x"74204e45",
  1763 => x"53000000",
  1764 => x"5363616e",
  1765 => x"6c696e65",
  1766 => x"73000000",
  1767 => x"48513258",
  1768 => x"2046696c",
  1769 => x"74657200",
  1770 => x"50312053",
  1771 => x"656c6563",
  1772 => x"74000000",
  1773 => x"50312053",
  1774 => x"74617274",
  1775 => x"00000000",
  1776 => x"4c6f6164",
  1777 => x"20524f4d",
  1778 => x"20100000",
  1779 => x"45786974",
  1780 => x"00000000",
  1781 => x"524f4d20",
  1782 => x"6c6f6164",
  1783 => x"696e6720",
  1784 => x"6661696c",
  1785 => x"65640000",
  1786 => x"4f4b0000",
  1787 => x"496e6974",
  1788 => x"69616c69",
  1789 => x"7a696e67",
  1790 => x"20534420",
  1791 => x"63617264",
  1792 => x"0a000000",
  1793 => x"16200000",
  1794 => x"14200000",
  1795 => x"15200000",
  1796 => x"53442069",
  1797 => x"6e69742e",
  1798 => x"2e2e0a00",
  1799 => x"53442063",
  1800 => x"61726420",
  1801 => x"72657365",
  1802 => x"74206661",
  1803 => x"696c6564",
  1804 => x"210a0000",
  1805 => x"53444843",
  1806 => x"20657272",
  1807 => x"6f72210a",
  1808 => x"00000000",
  1809 => x"57726974",
  1810 => x"65206661",
  1811 => x"696c6564",
  1812 => x"0a000000",
  1813 => x"52656164",
  1814 => x"20666169",
  1815 => x"6c65640a",
  1816 => x"00000000",
  1817 => x"43617264",
  1818 => x"20696e69",
  1819 => x"74206661",
  1820 => x"696c6564",
  1821 => x"0a000000",
  1822 => x"46415431",
  1823 => x"36202020",
  1824 => x"00000000",
  1825 => x"46415433",
  1826 => x"32202020",
  1827 => x"00000000",
  1828 => x"4e6f2070",
  1829 => x"61727469",
  1830 => x"74696f6e",
  1831 => x"20736967",
  1832 => x"0a000000",
  1833 => x"42616420",
  1834 => x"70617274",
  1835 => x"0a000000",
  1836 => x"4261636b",
  1837 => x"00000000",
  1838 => x"00000002",
  1839 => x"00000002",
  1840 => x"00001b84",
  1841 => x"0000034e",
  1842 => x"00000001",
  1843 => x"00001b90",
  1844 => x"00000000",
  1845 => x"00000001",
  1846 => x"00001b9c",
  1847 => x"00000001",
  1848 => x"00000002",
  1849 => x"00001ba8",
  1850 => x"00000362",
  1851 => x"00000002",
  1852 => x"00001bb4",
  1853 => x"00000373",
  1854 => x"00000002",
  1855 => x"00001bc0",
  1856 => x"00001b2e",
  1857 => x"00000002",
  1858 => x"00001bcc",
  1859 => x"00000774",
  1860 => x"00000000",
  1861 => x"00000000",
  1862 => x"00000000",
  1863 => x"00000004",
  1864 => x"00001bd4",
  1865 => x"00001d1c",
  1866 => x"00000004",
  1867 => x"00001be8",
  1868 => x"00001cbc",
  1869 => x"00000000",
  1870 => x"00000000",
  1871 => x"00000000",
  1872 => x"00000000",
  1873 => x"00000000",
  1874 => x"00000000",
  1875 => x"00000000",
  1876 => x"00000000",
  1877 => x"00000000",
  1878 => x"00000000",
  1879 => x"00000000",
  1880 => x"00000000",
  1881 => x"00000000",
  1882 => x"00000000",
  1883 => x"00000000",
  1884 => x"00000000",
  1885 => x"00000000",
  1886 => x"00000000",
  1887 => x"00000000",
  1888 => x"00000000",
  1889 => x"00000000",
  1890 => x"00000000",
  1891 => x"00000043",
  1892 => x"00000042",
  1893 => x"0000003b",
  1894 => x"0000004b",
  1895 => x"00000033",
  1896 => x"00000035",
  1897 => x"00000036",
  1898 => x"0000001e",
  1899 => x"0000001d",
  1900 => x"0000001b",
  1901 => x"0000001c",
  1902 => x"00000023",
  1903 => x"0000002b",
  1904 => x"0000002d",
  1905 => x"0000002e",
  1906 => x"00000016",
  1907 => x"00000000",
  1908 => x"00000000",
  1909 => x"00000002",
  1910 => x"0000223c",
  1911 => x"00001922",
  1912 => x"00000002",
  1913 => x"0000225a",
  1914 => x"00001922",
  1915 => x"00000002",
  1916 => x"00002278",
  1917 => x"00001922",
  1918 => x"00000002",
  1919 => x"00002296",
  1920 => x"00001922",
  1921 => x"00000002",
  1922 => x"000022b4",
  1923 => x"00001922",
  1924 => x"00000002",
  1925 => x"000022d2",
  1926 => x"00001922",
  1927 => x"00000002",
  1928 => x"000022f0",
  1929 => x"00001922",
  1930 => x"00000002",
  1931 => x"0000230e",
  1932 => x"00001922",
  1933 => x"00000002",
  1934 => x"0000232c",
  1935 => x"00001922",
  1936 => x"00000002",
  1937 => x"0000234a",
  1938 => x"00001922",
  1939 => x"00000002",
  1940 => x"00002368",
  1941 => x"00001922",
  1942 => x"00000002",
  1943 => x"00002386",
  1944 => x"00001922",
  1945 => x"00000002",
  1946 => x"000023a4",
  1947 => x"00001922",
  1948 => x"00000004",
  1949 => x"00001cb0",
  1950 => x"00000000",
  1951 => x"00000000",
  1952 => x"00000000",
  1953 => x"00001ac2",
  1954 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

