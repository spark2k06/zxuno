-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80d6",
     9 => x"94080b0b",
    10 => x"80d69808",
    11 => x"0b0b80d6",
    12 => x"9c080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"d69c0c0b",
    16 => x"0b80d698",
    17 => x"0c0b0b80",
    18 => x"d6940c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80cffc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80d69470",
    57 => x"80e0c827",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51a3cc",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80d6",
    65 => x"a40c9f0b",
    66 => x"80d6a80c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"d6a808ff",
    70 => x"0580d6a8",
    71 => x"0c80d6a8",
    72 => x"088025e8",
    73 => x"3880d6a4",
    74 => x"08ff0580",
    75 => x"d6a40c80",
    76 => x"d6a40880",
    77 => x"25d03880",
    78 => x"0b80d6a8",
    79 => x"0c800b80",
    80 => x"d6a40c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80d6a408",
   100 => x"25913882",
   101 => x"c82d80d6",
   102 => x"a408ff05",
   103 => x"80d6a40c",
   104 => x"838a0480",
   105 => x"d6a40880",
   106 => x"d6a80853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80d6a408",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"d6a80881",
   116 => x"0580d6a8",
   117 => x"0c80d6a8",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80d6a8",
   121 => x"0c80d6a4",
   122 => x"08810580",
   123 => x"d6a40c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480d6",
   128 => x"a8088105",
   129 => x"80d6a80c",
   130 => x"80d6a808",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80d6a8",
   134 => x"0c80d6a4",
   135 => x"08810580",
   136 => x"d6a40c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"d6ac0cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"d6ac0c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280d6",
   177 => x"ac088407",
   178 => x"80d6ac0c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80d2",
   183 => x"dc0c8171",
   184 => x"2bff05f6",
   185 => x"880cfecc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80d6ac",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80d6",
   208 => x"940c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"02dc050d",
  1093 => x"8059810b",
  1094 => x"ec0c840b",
  1095 => x"ec0c7a52",
  1096 => x"80d6b051",
  1097 => x"80c6cb2d",
  1098 => x"80d69408",
  1099 => x"792e80f4",
  1100 => x"3880d6b4",
  1101 => x"0879ff12",
  1102 => x"56595673",
  1103 => x"792e8b38",
  1104 => x"81187481",
  1105 => x"2a555873",
  1106 => x"f738f718",
  1107 => x"58815980",
  1108 => x"762580d0",
  1109 => x"38775273",
  1110 => x"5184a82d",
  1111 => x"80d78052",
  1112 => x"80d6b051",
  1113 => x"80c99f2d",
  1114 => x"80d69408",
  1115 => x"802e9b38",
  1116 => x"80d78057",
  1117 => x"83fc5576",
  1118 => x"70840558",
  1119 => x"08e80cfc",
  1120 => x"15557480",
  1121 => x"25f138a3",
  1122 => x"920480d6",
  1123 => x"94085984",
  1124 => x"805680d6",
  1125 => x"b05180c8",
  1126 => x"ee2dfc80",
  1127 => x"16811555",
  1128 => x"56a2cf04",
  1129 => x"80d6b408",
  1130 => x"f80c8051",
  1131 => x"86da2d78",
  1132 => x"802e8838",
  1133 => x"80d2e051",
  1134 => x"a3bf0480",
  1135 => x"d3e451ab",
  1136 => x"be2d7880",
  1137 => x"d6940c02",
  1138 => x"a4050d04",
  1139 => x"02f0050d",
  1140 => x"840bec0c",
  1141 => x"a8f02da5",
  1142 => x"a52d81f9",
  1143 => x"2d8352a8",
  1144 => x"d32d8151",
  1145 => x"858d2dff",
  1146 => x"12527180",
  1147 => x"25f13884",
  1148 => x"0bec0c80",
  1149 => x"d1905186",
  1150 => x"a02dbcfa",
  1151 => x"2d80d694",
  1152 => x"08802e81",
  1153 => x"8938a290",
  1154 => x"5180cff4",
  1155 => x"2d80d2e0",
  1156 => x"51abbe2d",
  1157 => x"a9922da5",
  1158 => x"b12dabd1",
  1159 => x"2d80d2f4",
  1160 => x"0b80f52d",
  1161 => x"80d4d008",
  1162 => x"70810654",
  1163 => x"55537180",
  1164 => x"2e853872",
  1165 => x"84075373",
  1166 => x"812a7081",
  1167 => x"06515271",
  1168 => x"802e8538",
  1169 => x"72820753",
  1170 => x"73822a70",
  1171 => x"81065152",
  1172 => x"71802e85",
  1173 => x"38728107",
  1174 => x"5373832a",
  1175 => x"70810651",
  1176 => x"5271802e",
  1177 => x"85387288",
  1178 => x"07537384",
  1179 => x"2a708106",
  1180 => x"51527180",
  1181 => x"2e853872",
  1182 => x"90075372",
  1183 => x"fc0c8652",
  1184 => x"80d69408",
  1185 => x"83388452",
  1186 => x"71ec0ca4",
  1187 => x"9704800b",
  1188 => x"80d6940c",
  1189 => x"0290050d",
  1190 => x"0471980c",
  1191 => x"04ffb008",
  1192 => x"80d6940c",
  1193 => x"04810bff",
  1194 => x"b00c0480",
  1195 => x"0bffb00c",
  1196 => x"0402f405",
  1197 => x"0da6bf04",
  1198 => x"80d69408",
  1199 => x"81f02e09",
  1200 => x"81068a38",
  1201 => x"810b80d4",
  1202 => x"c80ca6bf",
  1203 => x"0480d694",
  1204 => x"0881e02e",
  1205 => x"0981068a",
  1206 => x"38810b80",
  1207 => x"d4cc0ca6",
  1208 => x"bf0480d6",
  1209 => x"94085280",
  1210 => x"d4cc0880",
  1211 => x"2e893880",
  1212 => x"d6940881",
  1213 => x"80055271",
  1214 => x"842c728f",
  1215 => x"06535380",
  1216 => x"d4c80880",
  1217 => x"2e9a3872",
  1218 => x"842980d4",
  1219 => x"88057213",
  1220 => x"81712b70",
  1221 => x"09730806",
  1222 => x"730c5153",
  1223 => x"53a6b304",
  1224 => x"72842980",
  1225 => x"d4880572",
  1226 => x"1383712b",
  1227 => x"72080772",
  1228 => x"0c535380",
  1229 => x"0b80d4cc",
  1230 => x"0c800b80",
  1231 => x"d4c80c80",
  1232 => x"d6bc51a7",
  1233 => x"c62d80d6",
  1234 => x"9408ff24",
  1235 => x"feea3880",
  1236 => x"0b80d694",
  1237 => x"0c028c05",
  1238 => x"0d0402f8",
  1239 => x"050d80d4",
  1240 => x"88528f51",
  1241 => x"80727084",
  1242 => x"05540cff",
  1243 => x"11517080",
  1244 => x"25f23802",
  1245 => x"88050d04",
  1246 => x"02f0050d",
  1247 => x"7551a5ab",
  1248 => x"2d70822c",
  1249 => x"fc0680d4",
  1250 => x"88117210",
  1251 => x"9e067108",
  1252 => x"70722a70",
  1253 => x"83068274",
  1254 => x"2b700974",
  1255 => x"06760c54",
  1256 => x"51565753",
  1257 => x"5153a5a5",
  1258 => x"2d7180d6",
  1259 => x"940c0290",
  1260 => x"050d0402",
  1261 => x"fc050d72",
  1262 => x"5180710c",
  1263 => x"800b8412",
  1264 => x"0c028405",
  1265 => x"0d0402f0",
  1266 => x"050d7570",
  1267 => x"08841208",
  1268 => x"535353ff",
  1269 => x"5471712e",
  1270 => x"a838a5ab",
  1271 => x"2d841308",
  1272 => x"70842914",
  1273 => x"88117008",
  1274 => x"7081ff06",
  1275 => x"84180881",
  1276 => x"11870684",
  1277 => x"1a0c5351",
  1278 => x"55515151",
  1279 => x"a5a52d71",
  1280 => x"547380d6",
  1281 => x"940c0290",
  1282 => x"050d0402",
  1283 => x"f8050da5",
  1284 => x"ab2de008",
  1285 => x"708b2a70",
  1286 => x"81065152",
  1287 => x"5270802e",
  1288 => x"a13880d6",
  1289 => x"bc087084",
  1290 => x"2980d6c4",
  1291 => x"057381ff",
  1292 => x"06710c51",
  1293 => x"5180d6bc",
  1294 => x"08811187",
  1295 => x"0680d6bc",
  1296 => x"0c51800b",
  1297 => x"80d6e40c",
  1298 => x"a59d2da5",
  1299 => x"a52d0288",
  1300 => x"050d0402",
  1301 => x"fc050da5",
  1302 => x"ab2d810b",
  1303 => x"80d6e40c",
  1304 => x"a5a52d80",
  1305 => x"d6e40851",
  1306 => x"70f93802",
  1307 => x"84050d04",
  1308 => x"02fc050d",
  1309 => x"80d6bc51",
  1310 => x"a7b32da6",
  1311 => x"da2da88b",
  1312 => x"51a5992d",
  1313 => x"0284050d",
  1314 => x"0480d6ec",
  1315 => x"0880d694",
  1316 => x"0c0402fc",
  1317 => x"050d810b",
  1318 => x"80d4d40c",
  1319 => x"8151858d",
  1320 => x"2d028405",
  1321 => x"0d0402fc",
  1322 => x"050da9b0",
  1323 => x"04a5b12d",
  1324 => x"80f651a6",
  1325 => x"f82d80d6",
  1326 => x"9408f238",
  1327 => x"80da51a6",
  1328 => x"f82d80d6",
  1329 => x"9408e638",
  1330 => x"ab51a6f8",
  1331 => x"2d80d694",
  1332 => x"08db3880",
  1333 => x"d6940880",
  1334 => x"d4d40c80",
  1335 => x"d6940851",
  1336 => x"858d2d02",
  1337 => x"84050d04",
  1338 => x"02ec050d",
  1339 => x"76548052",
  1340 => x"870b8815",
  1341 => x"80f52d56",
  1342 => x"53747224",
  1343 => x"8338a053",
  1344 => x"72518384",
  1345 => x"2d81128b",
  1346 => x"1580f52d",
  1347 => x"54527272",
  1348 => x"25de3802",
  1349 => x"94050d04",
  1350 => x"02f0050d",
  1351 => x"80d6ec08",
  1352 => x"5481f92d",
  1353 => x"800b80d6",
  1354 => x"f00c7308",
  1355 => x"802e8189",
  1356 => x"38820b80",
  1357 => x"d6a80c80",
  1358 => x"d6f0088f",
  1359 => x"0680d6a4",
  1360 => x"0c730852",
  1361 => x"71832e96",
  1362 => x"38718326",
  1363 => x"89387181",
  1364 => x"2eb038ab",
  1365 => x"a2047185",
  1366 => x"2ea038ab",
  1367 => x"a2048814",
  1368 => x"80f52d84",
  1369 => x"150880d1",
  1370 => x"a8535452",
  1371 => x"86a02d71",
  1372 => x"84291370",
  1373 => x"085252ab",
  1374 => x"a6047351",
  1375 => x"a9e82dab",
  1376 => x"a20480d4",
  1377 => x"d0088815",
  1378 => x"082c7081",
  1379 => x"06515271",
  1380 => x"802e8838",
  1381 => x"80d1ac51",
  1382 => x"ab9f0480",
  1383 => x"d1b05186",
  1384 => x"a02d8414",
  1385 => x"085186a0",
  1386 => x"2d80d6f0",
  1387 => x"08810580",
  1388 => x"d6f00c8c",
  1389 => x"1454aaaa",
  1390 => x"04029005",
  1391 => x"0d047180",
  1392 => x"d6ec0caa",
  1393 => x"982d80d6",
  1394 => x"f008ff05",
  1395 => x"80d6f40c",
  1396 => x"0402e805",
  1397 => x"0d80d6ec",
  1398 => x"0880d6f8",
  1399 => x"08575580",
  1400 => x"f651a6f8",
  1401 => x"2d80d694",
  1402 => x"08812a70",
  1403 => x"81065152",
  1404 => x"71802ea4",
  1405 => x"38abfb04",
  1406 => x"a5b12d80",
  1407 => x"f651a6f8",
  1408 => x"2d80d694",
  1409 => x"08f23880",
  1410 => x"d4d40881",
  1411 => x"327080d4",
  1412 => x"d40c7052",
  1413 => x"52858d2d",
  1414 => x"800b80d6",
  1415 => x"e80c80d4",
  1416 => x"d40881f8",
  1417 => x"389d51a6",
  1418 => x"f82d80d6",
  1419 => x"9408802e",
  1420 => x"8b3880d6",
  1421 => x"e8088107",
  1422 => x"80d6e80c",
  1423 => x"9b51a6f8",
  1424 => x"2d80d694",
  1425 => x"08802e8b",
  1426 => x"3880d6e8",
  1427 => x"08820780",
  1428 => x"d6e80c9c",
  1429 => x"51a6f82d",
  1430 => x"80d69408",
  1431 => x"802e8b38",
  1432 => x"80d6e808",
  1433 => x"840780d6",
  1434 => x"e80ca351",
  1435 => x"a6f82d80",
  1436 => x"d6940880",
  1437 => x"2e8b3880",
  1438 => x"d6e80888",
  1439 => x"0780d6e8",
  1440 => x"0cab51a6",
  1441 => x"f82d80d6",
  1442 => x"9408802e",
  1443 => x"8b3880d6",
  1444 => x"e8089007",
  1445 => x"80d6e80c",
  1446 => x"80c351a6",
  1447 => x"f82d80d6",
  1448 => x"9408802e",
  1449 => x"8c3880d6",
  1450 => x"e8088280",
  1451 => x"0780d6e8",
  1452 => x"0c80c251",
  1453 => x"a6f82d80",
  1454 => x"d6940880",
  1455 => x"2e8c3880",
  1456 => x"d6e80884",
  1457 => x"800780d6",
  1458 => x"e80cbb51",
  1459 => x"a6f82d80",
  1460 => x"d6940880",
  1461 => x"2e8c3880",
  1462 => x"d6e80888",
  1463 => x"800780d6",
  1464 => x"e80c80cb",
  1465 => x"51a6f82d",
  1466 => x"80d69408",
  1467 => x"802e8c38",
  1468 => x"80d6e808",
  1469 => x"90800780",
  1470 => x"d6e80cb3",
  1471 => x"51a6f82d",
  1472 => x"80d69408",
  1473 => x"802e8c38",
  1474 => x"80d6e808",
  1475 => x"a0800780",
  1476 => x"d6e80c80",
  1477 => x"d6e808ed",
  1478 => x"0cb4d004",
  1479 => x"81f551a6",
  1480 => x"f82d80d6",
  1481 => x"9408812a",
  1482 => x"70810651",
  1483 => x"52719638",
  1484 => x"9d51a6f8",
  1485 => x"2d80d694",
  1486 => x"08812a70",
  1487 => x"81065152",
  1488 => x"71802eb3",
  1489 => x"3880d6f4",
  1490 => x"08527180",
  1491 => x"2e8a38ff",
  1492 => x"1280d6f4",
  1493 => x"0caef704",
  1494 => x"80d6f008",
  1495 => x"1080d6f0",
  1496 => x"08057084",
  1497 => x"29165152",
  1498 => x"88120880",
  1499 => x"2e8938ff",
  1500 => x"51881208",
  1501 => x"52712d81",
  1502 => x"f251a6f8",
  1503 => x"2d80d694",
  1504 => x"08812a70",
  1505 => x"81065152",
  1506 => x"7196389b",
  1507 => x"51a6f82d",
  1508 => x"80d69408",
  1509 => x"812a7081",
  1510 => x"06515271",
  1511 => x"802eb438",
  1512 => x"80d6f008",
  1513 => x"ff1180d6",
  1514 => x"f4085653",
  1515 => x"53737225",
  1516 => x"8a388114",
  1517 => x"80d6f40c",
  1518 => x"afd30472",
  1519 => x"10137084",
  1520 => x"29165152",
  1521 => x"88120880",
  1522 => x"2e8938fe",
  1523 => x"51881208",
  1524 => x"52712d81",
  1525 => x"fd51a6f8",
  1526 => x"2d80d694",
  1527 => x"08812a70",
  1528 => x"81065152",
  1529 => x"7196389c",
  1530 => x"51a6f82d",
  1531 => x"80d69408",
  1532 => x"812a7081",
  1533 => x"06515271",
  1534 => x"802eb138",
  1535 => x"80d6f408",
  1536 => x"802e8a38",
  1537 => x"800b80d6",
  1538 => x"f40cb0ac",
  1539 => x"0480d6f0",
  1540 => x"081080d6",
  1541 => x"f0080570",
  1542 => x"84291651",
  1543 => x"52881208",
  1544 => x"802e8938",
  1545 => x"fd518812",
  1546 => x"0852712d",
  1547 => x"81fa51a6",
  1548 => x"f82d80d6",
  1549 => x"9408812a",
  1550 => x"70810651",
  1551 => x"52719638",
  1552 => x"a351a6f8",
  1553 => x"2d80d694",
  1554 => x"08812a70",
  1555 => x"81065152",
  1556 => x"71802eb1",
  1557 => x"3880d6f0",
  1558 => x"08ff1154",
  1559 => x"5280d6f4",
  1560 => x"08732589",
  1561 => x"387280d6",
  1562 => x"f40cb185",
  1563 => x"04711012",
  1564 => x"70842916",
  1565 => x"51528812",
  1566 => x"08802e89",
  1567 => x"38fc5188",
  1568 => x"12085271",
  1569 => x"2d80d6f4",
  1570 => x"08705354",
  1571 => x"73802e8a",
  1572 => x"388c15ff",
  1573 => x"155555b1",
  1574 => x"8c04820b",
  1575 => x"80d6a80c",
  1576 => x"718f0680",
  1577 => x"d6a40c81",
  1578 => x"eb51a6f8",
  1579 => x"2d80d694",
  1580 => x"08812a70",
  1581 => x"81065152",
  1582 => x"71802ead",
  1583 => x"38740885",
  1584 => x"2e098106",
  1585 => x"a4388815",
  1586 => x"80f52dff",
  1587 => x"05527188",
  1588 => x"1681b72d",
  1589 => x"71982b52",
  1590 => x"71802588",
  1591 => x"38800b88",
  1592 => x"1681b72d",
  1593 => x"7451a9e8",
  1594 => x"2d81f451",
  1595 => x"a6f82d80",
  1596 => x"d6940881",
  1597 => x"2a708106",
  1598 => x"51527180",
  1599 => x"2eb33874",
  1600 => x"08852e09",
  1601 => x"8106aa38",
  1602 => x"881580f5",
  1603 => x"2d810552",
  1604 => x"71881681",
  1605 => x"b72d7181",
  1606 => x"ff068b16",
  1607 => x"80f52d54",
  1608 => x"52727227",
  1609 => x"87387288",
  1610 => x"1681b72d",
  1611 => x"7451a9e8",
  1612 => x"2d80da51",
  1613 => x"a6f82d80",
  1614 => x"d6940881",
  1615 => x"2a708106",
  1616 => x"51527197",
  1617 => x"38ab51a6",
  1618 => x"f82d80d6",
  1619 => x"9408812a",
  1620 => x"70810651",
  1621 => x"5271802e",
  1622 => x"81ad3880",
  1623 => x"d6ec0880",
  1624 => x"d6f40855",
  1625 => x"5373802e",
  1626 => x"8a388c13",
  1627 => x"ff155553",
  1628 => x"b2e50472",
  1629 => x"08527182",
  1630 => x"2ea63871",
  1631 => x"82268938",
  1632 => x"71812eaa",
  1633 => x"38b48704",
  1634 => x"71832eb4",
  1635 => x"3871842e",
  1636 => x"09810680",
  1637 => x"f2388813",
  1638 => x"0851abbe",
  1639 => x"2db48704",
  1640 => x"80d6f408",
  1641 => x"51881308",
  1642 => x"52712db4",
  1643 => x"8704810b",
  1644 => x"8814082b",
  1645 => x"80d4d008",
  1646 => x"3280d4d0",
  1647 => x"0cb3db04",
  1648 => x"881380f5",
  1649 => x"2d81058b",
  1650 => x"1480f52d",
  1651 => x"53547174",
  1652 => x"24833880",
  1653 => x"54738814",
  1654 => x"81b72daa",
  1655 => x"982db487",
  1656 => x"04750880",
  1657 => x"2ea43875",
  1658 => x"0851a6f8",
  1659 => x"2d80d694",
  1660 => x"08810652",
  1661 => x"71802e8c",
  1662 => x"3880d6f4",
  1663 => x"08518416",
  1664 => x"0852712d",
  1665 => x"88165675",
  1666 => x"d8388054",
  1667 => x"800b80d6",
  1668 => x"a80c738f",
  1669 => x"0680d6a4",
  1670 => x"0ca05273",
  1671 => x"80d6f408",
  1672 => x"2e098106",
  1673 => x"993880d6",
  1674 => x"f008ff05",
  1675 => x"74327009",
  1676 => x"81057072",
  1677 => x"079f2a91",
  1678 => x"71315151",
  1679 => x"53537151",
  1680 => x"83842d81",
  1681 => x"14548e74",
  1682 => x"25c23880",
  1683 => x"d4d40852",
  1684 => x"7180d694",
  1685 => x"0c029805",
  1686 => x"0d0402f4",
  1687 => x"050dd452",
  1688 => x"81ff720c",
  1689 => x"71085381",
  1690 => x"ff720c72",
  1691 => x"882b83fe",
  1692 => x"80067208",
  1693 => x"7081ff06",
  1694 => x"51525381",
  1695 => x"ff720c72",
  1696 => x"7107882b",
  1697 => x"72087081",
  1698 => x"ff065152",
  1699 => x"5381ff72",
  1700 => x"0c727107",
  1701 => x"882b7208",
  1702 => x"7081ff06",
  1703 => x"720780d6",
  1704 => x"940c5253",
  1705 => x"028c050d",
  1706 => x"0402f405",
  1707 => x"0d747671",
  1708 => x"81ff06d4",
  1709 => x"0c535380",
  1710 => x"d6fc0885",
  1711 => x"3871892b",
  1712 => x"5271982a",
  1713 => x"d40c7190",
  1714 => x"2a7081ff",
  1715 => x"06d40c51",
  1716 => x"71882a70",
  1717 => x"81ff06d4",
  1718 => x"0c517181",
  1719 => x"ff06d40c",
  1720 => x"72902a70",
  1721 => x"81ff06d4",
  1722 => x"0c51d408",
  1723 => x"7081ff06",
  1724 => x"515182b8",
  1725 => x"bf527081",
  1726 => x"ff2e0981",
  1727 => x"06943881",
  1728 => x"ff0bd40c",
  1729 => x"d4087081",
  1730 => x"ff06ff14",
  1731 => x"54515171",
  1732 => x"e5387080",
  1733 => x"d6940c02",
  1734 => x"8c050d04",
  1735 => x"02fc050d",
  1736 => x"81c75181",
  1737 => x"ff0bd40c",
  1738 => x"ff115170",
  1739 => x"8025f438",
  1740 => x"0284050d",
  1741 => x"0402f405",
  1742 => x"0d81ff0b",
  1743 => x"d40c9353",
  1744 => x"805287fc",
  1745 => x"80c151b5",
  1746 => x"a92d80d6",
  1747 => x"94088b38",
  1748 => x"81ff0bd4",
  1749 => x"0c8153b6",
  1750 => x"e304b69c",
  1751 => x"2dff1353",
  1752 => x"72de3872",
  1753 => x"80d6940c",
  1754 => x"028c050d",
  1755 => x"0402ec05",
  1756 => x"0d810b80",
  1757 => x"d6fc0c84",
  1758 => x"54d00870",
  1759 => x"8f2a7081",
  1760 => x"06515153",
  1761 => x"72f33872",
  1762 => x"d00cb69c",
  1763 => x"2d80d1b4",
  1764 => x"5186a02d",
  1765 => x"d008708f",
  1766 => x"2a708106",
  1767 => x"51515372",
  1768 => x"f338810b",
  1769 => x"d00cb153",
  1770 => x"805284d4",
  1771 => x"80c051b5",
  1772 => x"a92d80d6",
  1773 => x"9408812e",
  1774 => x"93387282",
  1775 => x"2ebf38ff",
  1776 => x"135372e4",
  1777 => x"38ff1454",
  1778 => x"73ffae38",
  1779 => x"b69c2d83",
  1780 => x"aa52849c",
  1781 => x"80c851b5",
  1782 => x"a92d80d6",
  1783 => x"9408812e",
  1784 => x"09810693",
  1785 => x"38b4da2d",
  1786 => x"80d69408",
  1787 => x"83ffff06",
  1788 => x"537283aa",
  1789 => x"2e9f38b6",
  1790 => x"b52db890",
  1791 => x"0480d1c0",
  1792 => x"5186a02d",
  1793 => x"8053b9e5",
  1794 => x"0480d1d8",
  1795 => x"5186a02d",
  1796 => x"8054b9b6",
  1797 => x"0481ff0b",
  1798 => x"d40cb154",
  1799 => x"b69c2d8f",
  1800 => x"cf538052",
  1801 => x"87fc80f7",
  1802 => x"51b5a92d",
  1803 => x"80d69408",
  1804 => x"5580d694",
  1805 => x"08812e09",
  1806 => x"81069c38",
  1807 => x"81ff0bd4",
  1808 => x"0c820a52",
  1809 => x"849c80e9",
  1810 => x"51b5a92d",
  1811 => x"80d69408",
  1812 => x"802e8d38",
  1813 => x"b69c2dff",
  1814 => x"135372c6",
  1815 => x"38b9a904",
  1816 => x"81ff0bd4",
  1817 => x"0c80d694",
  1818 => x"085287fc",
  1819 => x"80fa51b5",
  1820 => x"a92d80d6",
  1821 => x"9408b238",
  1822 => x"81ff0bd4",
  1823 => x"0cd40853",
  1824 => x"81ff0bd4",
  1825 => x"0c81ff0b",
  1826 => x"d40c81ff",
  1827 => x"0bd40c81",
  1828 => x"ff0bd40c",
  1829 => x"72862a70",
  1830 => x"81067656",
  1831 => x"51537296",
  1832 => x"3880d694",
  1833 => x"0854b9b6",
  1834 => x"0473822e",
  1835 => x"fedb38ff",
  1836 => x"145473fe",
  1837 => x"e7387380",
  1838 => x"d6fc0c73",
  1839 => x"8b388152",
  1840 => x"87fc80d0",
  1841 => x"51b5a92d",
  1842 => x"81ff0bd4",
  1843 => x"0cd00870",
  1844 => x"8f2a7081",
  1845 => x"06515153",
  1846 => x"72f33872",
  1847 => x"d00c81ff",
  1848 => x"0bd40c81",
  1849 => x"537280d6",
  1850 => x"940c0294",
  1851 => x"050d0402",
  1852 => x"e8050d78",
  1853 => x"55805681",
  1854 => x"ff0bd40c",
  1855 => x"d008708f",
  1856 => x"2a708106",
  1857 => x"51515372",
  1858 => x"f3388281",
  1859 => x"0bd00c81",
  1860 => x"ff0bd40c",
  1861 => x"775287fc",
  1862 => x"80d151b5",
  1863 => x"a92d80db",
  1864 => x"c6df5480",
  1865 => x"d6940880",
  1866 => x"2e8b3880",
  1867 => x"d1f85186",
  1868 => x"a02dbb89",
  1869 => x"0481ff0b",
  1870 => x"d40cd408",
  1871 => x"7081ff06",
  1872 => x"51537281",
  1873 => x"fe2e0981",
  1874 => x"069e3880",
  1875 => x"ff53b4da",
  1876 => x"2d80d694",
  1877 => x"08757084",
  1878 => x"05570cff",
  1879 => x"13537280",
  1880 => x"25ec3881",
  1881 => x"56baee04",
  1882 => x"ff145473",
  1883 => x"c83881ff",
  1884 => x"0bd40c81",
  1885 => x"ff0bd40c",
  1886 => x"d008708f",
  1887 => x"2a708106",
  1888 => x"51515372",
  1889 => x"f33872d0",
  1890 => x"0c7580d6",
  1891 => x"940c0298",
  1892 => x"050d0402",
  1893 => x"e8050d77",
  1894 => x"797b5855",
  1895 => x"55805372",
  1896 => x"7625a338",
  1897 => x"74708105",
  1898 => x"5680f52d",
  1899 => x"74708105",
  1900 => x"5680f52d",
  1901 => x"52527171",
  1902 => x"2e863881",
  1903 => x"51bbc804",
  1904 => x"811353bb",
  1905 => x"9f048051",
  1906 => x"7080d694",
  1907 => x"0c029805",
  1908 => x"0d0402ec",
  1909 => x"050d7655",
  1910 => x"74802e80",
  1911 => x"c4389a15",
  1912 => x"80e02d51",
  1913 => x"80c9f92d",
  1914 => x"80d69408",
  1915 => x"80d69408",
  1916 => x"80ddb00c",
  1917 => x"80d69408",
  1918 => x"545480dd",
  1919 => x"8c08802e",
  1920 => x"9b389415",
  1921 => x"80e02d51",
  1922 => x"80c9f92d",
  1923 => x"80d69408",
  1924 => x"902b83ff",
  1925 => x"f00a0670",
  1926 => x"75075153",
  1927 => x"7280ddb0",
  1928 => x"0c80ddb0",
  1929 => x"08537280",
  1930 => x"2e9d3880",
  1931 => x"dd8408fe",
  1932 => x"14712980",
  1933 => x"dd980805",
  1934 => x"80ddb40c",
  1935 => x"70842b80",
  1936 => x"dd900c54",
  1937 => x"bcf50480",
  1938 => x"dd9c0880",
  1939 => x"ddb00c80",
  1940 => x"dda00880",
  1941 => x"ddb40c80",
  1942 => x"dd8c0880",
  1943 => x"2e8b3880",
  1944 => x"dd840884",
  1945 => x"2b53bcf0",
  1946 => x"0480dda4",
  1947 => x"08842b53",
  1948 => x"7280dd90",
  1949 => x"0c029405",
  1950 => x"0d0402d8",
  1951 => x"050d800b",
  1952 => x"80dd8c0c",
  1953 => x"8454b6ed",
  1954 => x"2d80d694",
  1955 => x"08802e97",
  1956 => x"3880d780",
  1957 => x"528051b9",
  1958 => x"ef2d80d6",
  1959 => x"9408802e",
  1960 => x"8638fe54",
  1961 => x"bdaf04ff",
  1962 => x"14547380",
  1963 => x"24d83873",
  1964 => x"8e3880d2",
  1965 => x"885186a0",
  1966 => x"2d735580",
  1967 => x"c3890480",
  1968 => x"56810b80",
  1969 => x"ddb80c88",
  1970 => x"5380d29c",
  1971 => x"5280d7b6",
  1972 => x"51bb932d",
  1973 => x"80d69408",
  1974 => x"762e0981",
  1975 => x"06893880",
  1976 => x"d6940880",
  1977 => x"ddb80c88",
  1978 => x"5380d2a8",
  1979 => x"5280d7d2",
  1980 => x"51bb932d",
  1981 => x"80d69408",
  1982 => x"893880d6",
  1983 => x"940880dd",
  1984 => x"b80c80dd",
  1985 => x"b808802e",
  1986 => x"81823880",
  1987 => x"dac60b80",
  1988 => x"f52d80da",
  1989 => x"c70b80f5",
  1990 => x"2d71982b",
  1991 => x"71902b07",
  1992 => x"80dac80b",
  1993 => x"80f52d70",
  1994 => x"882b7207",
  1995 => x"80dac90b",
  1996 => x"80f52d71",
  1997 => x"0780dafe",
  1998 => x"0b80f52d",
  1999 => x"80daff0b",
  2000 => x"80f52d71",
  2001 => x"882b0753",
  2002 => x"5f54525a",
  2003 => x"56575573",
  2004 => x"81abaa2e",
  2005 => x"0981068f",
  2006 => x"38755180",
  2007 => x"c9c82d80",
  2008 => x"d6940856",
  2009 => x"bef50473",
  2010 => x"82d4d52e",
  2011 => x"883880d2",
  2012 => x"b451bfc1",
  2013 => x"0480d780",
  2014 => x"527551b9",
  2015 => x"ef2d80d6",
  2016 => x"94085580",
  2017 => x"d6940880",
  2018 => x"2e83fe38",
  2019 => x"885380d2",
  2020 => x"a85280d7",
  2021 => x"d251bb93",
  2022 => x"2d80d694",
  2023 => x"088a3881",
  2024 => x"0b80dd8c",
  2025 => x"0cbfc804",
  2026 => x"885380d2",
  2027 => x"9c5280d7",
  2028 => x"b651bb93",
  2029 => x"2d80d694",
  2030 => x"08802e8c",
  2031 => x"3880d2c8",
  2032 => x"5186a02d",
  2033 => x"80c0a704",
  2034 => x"80dafe0b",
  2035 => x"80f52d54",
  2036 => x"7380d52e",
  2037 => x"09810680",
  2038 => x"ce3880da",
  2039 => x"ff0b80f5",
  2040 => x"2d547381",
  2041 => x"aa2e0981",
  2042 => x"06bd3880",
  2043 => x"0b80d780",
  2044 => x"0b80f52d",
  2045 => x"56547481",
  2046 => x"e92e8338",
  2047 => x"81547481",
  2048 => x"eb2e8c38",
  2049 => x"80557375",
  2050 => x"2e098106",
  2051 => x"82fb3880",
  2052 => x"d78b0b80",
  2053 => x"f52d5574",
  2054 => x"8e3880d7",
  2055 => x"8c0b80f5",
  2056 => x"2d547382",
  2057 => x"2e873880",
  2058 => x"5580c389",
  2059 => x"0480d78d",
  2060 => x"0b80f52d",
  2061 => x"7080dd84",
  2062 => x"0cff0580",
  2063 => x"dd880c80",
  2064 => x"d78e0b80",
  2065 => x"f52d80d7",
  2066 => x"8f0b80f5",
  2067 => x"2d587605",
  2068 => x"77828029",
  2069 => x"057080dd",
  2070 => x"940c80d7",
  2071 => x"900b80f5",
  2072 => x"2d7080dd",
  2073 => x"a80c80dd",
  2074 => x"8c085957",
  2075 => x"5876802e",
  2076 => x"81b83888",
  2077 => x"5380d2a8",
  2078 => x"5280d7d2",
  2079 => x"51bb932d",
  2080 => x"80d69408",
  2081 => x"82833880",
  2082 => x"dd840870",
  2083 => x"842b80dd",
  2084 => x"900c7080",
  2085 => x"dda40c80",
  2086 => x"d7a50b80",
  2087 => x"f52d80d7",
  2088 => x"a40b80f5",
  2089 => x"2d718280",
  2090 => x"290580d7",
  2091 => x"a60b80f5",
  2092 => x"2d708480",
  2093 => x"80291280",
  2094 => x"d7a70b80",
  2095 => x"f52d7081",
  2096 => x"800a2912",
  2097 => x"7080ddac",
  2098 => x"0c80dda8",
  2099 => x"08712980",
  2100 => x"dd940805",
  2101 => x"7080dd98",
  2102 => x"0c80d7ad",
  2103 => x"0b80f52d",
  2104 => x"80d7ac0b",
  2105 => x"80f52d71",
  2106 => x"82802905",
  2107 => x"80d7ae0b",
  2108 => x"80f52d70",
  2109 => x"84808029",
  2110 => x"1280d7af",
  2111 => x"0b80f52d",
  2112 => x"70982b81",
  2113 => x"f00a0672",
  2114 => x"057080dd",
  2115 => x"9c0cfe11",
  2116 => x"7e297705",
  2117 => x"80dda00c",
  2118 => x"52595243",
  2119 => x"545e5152",
  2120 => x"59525d57",
  2121 => x"595780c3",
  2122 => x"820480d7",
  2123 => x"920b80f5",
  2124 => x"2d80d791",
  2125 => x"0b80f52d",
  2126 => x"71828029",
  2127 => x"057080dd",
  2128 => x"900c70a0",
  2129 => x"2983ff05",
  2130 => x"70892a70",
  2131 => x"80dda40c",
  2132 => x"80d7970b",
  2133 => x"80f52d80",
  2134 => x"d7960b80",
  2135 => x"f52d7182",
  2136 => x"80290570",
  2137 => x"80ddac0c",
  2138 => x"7b71291e",
  2139 => x"7080dda0",
  2140 => x"0c7d80dd",
  2141 => x"9c0c7305",
  2142 => x"80dd980c",
  2143 => x"555e5151",
  2144 => x"55558051",
  2145 => x"bbd22d81",
  2146 => x"557480d6",
  2147 => x"940c02a8",
  2148 => x"050d0402",
  2149 => x"ec050d76",
  2150 => x"70872c71",
  2151 => x"80ff0655",
  2152 => x"565480dd",
  2153 => x"8c088a38",
  2154 => x"73882c74",
  2155 => x"81ff0654",
  2156 => x"5580d780",
  2157 => x"5280dd94",
  2158 => x"081551b9",
  2159 => x"ef2d80d6",
  2160 => x"94085480",
  2161 => x"d6940880",
  2162 => x"2ebb3880",
  2163 => x"dd8c0880",
  2164 => x"2e9c3872",
  2165 => x"842980d7",
  2166 => x"80057008",
  2167 => x"525380c9",
  2168 => x"c82d80d6",
  2169 => x"9408f00a",
  2170 => x"065380c4",
  2171 => x"83047210",
  2172 => x"80d78005",
  2173 => x"7080e02d",
  2174 => x"525380c9",
  2175 => x"f92d80d6",
  2176 => x"94085372",
  2177 => x"547380d6",
  2178 => x"940c0294",
  2179 => x"050d0402",
  2180 => x"e0050d79",
  2181 => x"70842c80",
  2182 => x"ddb40805",
  2183 => x"718f0652",
  2184 => x"5553728a",
  2185 => x"3880d780",
  2186 => x"527351b9",
  2187 => x"ef2d72a0",
  2188 => x"2980d780",
  2189 => x"05548074",
  2190 => x"80f52d56",
  2191 => x"5374732e",
  2192 => x"83388153",
  2193 => x"7481e52e",
  2194 => x"81f53881",
  2195 => x"70740654",
  2196 => x"5872802e",
  2197 => x"81e9388b",
  2198 => x"1480f52d",
  2199 => x"70832a79",
  2200 => x"06585676",
  2201 => x"9c3880d4",
  2202 => x"d8085372",
  2203 => x"89387280",
  2204 => x"db800b81",
  2205 => x"b72d7680",
  2206 => x"d4d80c73",
  2207 => x"5380c6c1",
  2208 => x"04758f2e",
  2209 => x"09810681",
  2210 => x"b638749f",
  2211 => x"068d2980",
  2212 => x"daf31151",
  2213 => x"53811480",
  2214 => x"f52d7370",
  2215 => x"81055581",
  2216 => x"b72d8314",
  2217 => x"80f52d73",
  2218 => x"70810555",
  2219 => x"81b72d85",
  2220 => x"1480f52d",
  2221 => x"73708105",
  2222 => x"5581b72d",
  2223 => x"871480f5",
  2224 => x"2d737081",
  2225 => x"055581b7",
  2226 => x"2d891480",
  2227 => x"f52d7370",
  2228 => x"81055581",
  2229 => x"b72d8e14",
  2230 => x"80f52d73",
  2231 => x"70810555",
  2232 => x"81b72d90",
  2233 => x"1480f52d",
  2234 => x"73708105",
  2235 => x"5581b72d",
  2236 => x"921480f5",
  2237 => x"2d737081",
  2238 => x"055581b7",
  2239 => x"2d941480",
  2240 => x"f52d7370",
  2241 => x"81055581",
  2242 => x"b72d9614",
  2243 => x"80f52d73",
  2244 => x"70810555",
  2245 => x"81b72d98",
  2246 => x"1480f52d",
  2247 => x"73708105",
  2248 => x"5581b72d",
  2249 => x"9c1480f5",
  2250 => x"2d737081",
  2251 => x"055581b7",
  2252 => x"2d9e1480",
  2253 => x"f52d7381",
  2254 => x"b72d7780",
  2255 => x"d4d80c80",
  2256 => x"537280d6",
  2257 => x"940c02a0",
  2258 => x"050d0402",
  2259 => x"cc050d7e",
  2260 => x"605e5a80",
  2261 => x"0b80ddb0",
  2262 => x"0880ddb4",
  2263 => x"08595c56",
  2264 => x"805880dd",
  2265 => x"9008782e",
  2266 => x"81bc3877",
  2267 => x"8f06a017",
  2268 => x"57547391",
  2269 => x"3880d780",
  2270 => x"52765181",
  2271 => x"1757b9ef",
  2272 => x"2d80d780",
  2273 => x"56807680",
  2274 => x"f52d5654",
  2275 => x"74742e83",
  2276 => x"38815474",
  2277 => x"81e52e81",
  2278 => x"81388170",
  2279 => x"7506555c",
  2280 => x"73802e80",
  2281 => x"f5388b16",
  2282 => x"80f52d98",
  2283 => x"06597880",
  2284 => x"e9388b53",
  2285 => x"7c527551",
  2286 => x"bb932d80",
  2287 => x"d6940880",
  2288 => x"d9389c16",
  2289 => x"085180c9",
  2290 => x"c82d80d6",
  2291 => x"9408841b",
  2292 => x"0c9a1680",
  2293 => x"e02d5180",
  2294 => x"c9f92d80",
  2295 => x"d6940880",
  2296 => x"d6940888",
  2297 => x"1c0c80d6",
  2298 => x"94085555",
  2299 => x"80dd8c08",
  2300 => x"802e9a38",
  2301 => x"941680e0",
  2302 => x"2d5180c9",
  2303 => x"f92d80d6",
  2304 => x"9408902b",
  2305 => x"83fff00a",
  2306 => x"06701651",
  2307 => x"5473881b",
  2308 => x"0c787a0c",
  2309 => x"7b5480c8",
  2310 => x"e4048118",
  2311 => x"5880dd90",
  2312 => x"087826fe",
  2313 => x"c63880dd",
  2314 => x"8c08802e",
  2315 => x"b5387a51",
  2316 => x"80c3932d",
  2317 => x"80d69408",
  2318 => x"80d69408",
  2319 => x"80ffffff",
  2320 => x"f806555b",
  2321 => x"7380ffff",
  2322 => x"fff82e96",
  2323 => x"3880d694",
  2324 => x"08fe0580",
  2325 => x"dd840829",
  2326 => x"80dd9808",
  2327 => x"055780c6",
  2328 => x"e0048054",
  2329 => x"7380d694",
  2330 => x"0c02b405",
  2331 => x"0d0402f4",
  2332 => x"050d7470",
  2333 => x"08810571",
  2334 => x"0c700880",
  2335 => x"dd880806",
  2336 => x"53537190",
  2337 => x"38881308",
  2338 => x"5180c393",
  2339 => x"2d80d694",
  2340 => x"0888140c",
  2341 => x"810b80d6",
  2342 => x"940c028c",
  2343 => x"050d0402",
  2344 => x"f0050d75",
  2345 => x"881108fe",
  2346 => x"0580dd84",
  2347 => x"082980dd",
  2348 => x"98081172",
  2349 => x"0880dd88",
  2350 => x"08060579",
  2351 => x"55535454",
  2352 => x"b9ef2d02",
  2353 => x"90050d04",
  2354 => x"02f4050d",
  2355 => x"7470882a",
  2356 => x"83fe8006",
  2357 => x"7072982a",
  2358 => x"0772882b",
  2359 => x"87fc8080",
  2360 => x"0673982b",
  2361 => x"81f00a06",
  2362 => x"71730707",
  2363 => x"80d6940c",
  2364 => x"56515351",
  2365 => x"028c050d",
  2366 => x"0402f805",
  2367 => x"0d028e05",
  2368 => x"80f52d74",
  2369 => x"882b0770",
  2370 => x"83ffff06",
  2371 => x"80d6940c",
  2372 => x"51028805",
  2373 => x"0d0402f4",
  2374 => x"050d7476",
  2375 => x"78535452",
  2376 => x"80712597",
  2377 => x"38727081",
  2378 => x"055480f5",
  2379 => x"2d727081",
  2380 => x"055481b7",
  2381 => x"2dff1151",
  2382 => x"70eb3880",
  2383 => x"7281b72d",
  2384 => x"028c050d",
  2385 => x"0402e805",
  2386 => x"0d775680",
  2387 => x"70565473",
  2388 => x"7624b738",
  2389 => x"80dd9008",
  2390 => x"742eaf38",
  2391 => x"735180c4",
  2392 => x"8f2d80d6",
  2393 => x"940880d6",
  2394 => x"94080981",
  2395 => x"057080d6",
  2396 => x"9408079f",
  2397 => x"2a770581",
  2398 => x"17575753",
  2399 => x"53747624",
  2400 => x"893880dd",
  2401 => x"90087426",
  2402 => x"d3387280",
  2403 => x"d6940c02",
  2404 => x"98050d04",
  2405 => x"02f0050d",
  2406 => x"80d69008",
  2407 => x"165180ca",
  2408 => x"c52d80d6",
  2409 => x"9408802e",
  2410 => x"a0388b53",
  2411 => x"80d69408",
  2412 => x"5280db80",
  2413 => x"5180ca96",
  2414 => x"2d80ddbc",
  2415 => x"08547380",
  2416 => x"2e873880",
  2417 => x"db805173",
  2418 => x"2d029005",
  2419 => x"0d0402dc",
  2420 => x"050d8070",
  2421 => x"5a557480",
  2422 => x"d6900825",
  2423 => x"b53880dd",
  2424 => x"9008752e",
  2425 => x"ad387851",
  2426 => x"80c48f2d",
  2427 => x"80d69408",
  2428 => x"09810570",
  2429 => x"80d69408",
  2430 => x"079f2a76",
  2431 => x"05811b5b",
  2432 => x"56547480",
  2433 => x"d6900825",
  2434 => x"893880dd",
  2435 => x"90087926",
  2436 => x"d5388055",
  2437 => x"7880dd90",
  2438 => x"082781e4",
  2439 => x"38785180",
  2440 => x"c48f2d80",
  2441 => x"d6940880",
  2442 => x"2e81b438",
  2443 => x"80d69408",
  2444 => x"8b0580f5",
  2445 => x"2d70842a",
  2446 => x"70810677",
  2447 => x"1078842b",
  2448 => x"80db800b",
  2449 => x"80f52d5c",
  2450 => x"5c535155",
  2451 => x"5673802e",
  2452 => x"80ce3874",
  2453 => x"16822b80",
  2454 => x"cea40b80",
  2455 => x"d4e4120c",
  2456 => x"54777531",
  2457 => x"1080ddc0",
  2458 => x"11555690",
  2459 => x"74708105",
  2460 => x"5681b72d",
  2461 => x"a07481b7",
  2462 => x"2d7681ff",
  2463 => x"06811658",
  2464 => x"5473802e",
  2465 => x"8b389c53",
  2466 => x"80db8052",
  2467 => x"80cd9704",
  2468 => x"8b5380d6",
  2469 => x"94085280",
  2470 => x"ddc21651",
  2471 => x"80cdd504",
  2472 => x"7416822b",
  2473 => x"80cb940b",
  2474 => x"80d4e412",
  2475 => x"0c547681",
  2476 => x"ff068116",
  2477 => x"58547380",
  2478 => x"2e8b389c",
  2479 => x"5380db80",
  2480 => x"5280cdcc",
  2481 => x"048b5380",
  2482 => x"d6940852",
  2483 => x"77753110",
  2484 => x"80ddc005",
  2485 => x"51765580",
  2486 => x"ca962d80",
  2487 => x"cdf40474",
  2488 => x"90297531",
  2489 => x"701080dd",
  2490 => x"c0055154",
  2491 => x"80d69408",
  2492 => x"7481b72d",
  2493 => x"81195974",
  2494 => x"8b24a438",
  2495 => x"80cc9404",
  2496 => x"74902975",
  2497 => x"31701080",
  2498 => x"ddc0058c",
  2499 => x"77315751",
  2500 => x"54807481",
  2501 => x"b72d9e14",
  2502 => x"ff165654",
  2503 => x"74f33802",
  2504 => x"a4050d04",
  2505 => x"02fc050d",
  2506 => x"80d69008",
  2507 => x"135180ca",
  2508 => x"c52d80d6",
  2509 => x"9408802e",
  2510 => x"893880d6",
  2511 => x"940851bb",
  2512 => x"d22d800b",
  2513 => x"80d6900c",
  2514 => x"80cbce2d",
  2515 => x"aa982d02",
  2516 => x"84050d04",
  2517 => x"02fc050d",
  2518 => x"725170fd",
  2519 => x"2eb23870",
  2520 => x"fd248b38",
  2521 => x"70fc2e80",
  2522 => x"d03880cf",
  2523 => x"c30470fe",
  2524 => x"2eb93870",
  2525 => x"ff2e0981",
  2526 => x"0680c838",
  2527 => x"80d69008",
  2528 => x"5170802e",
  2529 => x"be38ff11",
  2530 => x"80d6900c",
  2531 => x"80cfc304",
  2532 => x"80d69008",
  2533 => x"f0057080",
  2534 => x"d6900c51",
  2535 => x"708025a3",
  2536 => x"38800b80",
  2537 => x"d6900c80",
  2538 => x"cfc30480",
  2539 => x"d6900881",
  2540 => x"0580d690",
  2541 => x"0c80cfc3",
  2542 => x"0480d690",
  2543 => x"08900580",
  2544 => x"d6900c80",
  2545 => x"cbce2daa",
  2546 => x"982d0284",
  2547 => x"050d0402",
  2548 => x"fc050d80",
  2549 => x"0b80d690",
  2550 => x"0c80cbce",
  2551 => x"2da9892d",
  2552 => x"80d69408",
  2553 => x"80d6800c",
  2554 => x"80d4dc51",
  2555 => x"abbe2d02",
  2556 => x"84050d04",
  2557 => x"7180ddbc",
  2558 => x"0c040000",
  2559 => x"00ffffff",
  2560 => x"ff00ffff",
  2561 => x"ffff00ff",
  2562 => x"ffffff00",
  2563 => x"52657365",
  2564 => x"74000000",
  2565 => x"5363616e",
  2566 => x"6c696e65",
  2567 => x"73000000",
  2568 => x"50414c20",
  2569 => x"2f204e54",
  2570 => x"53430000",
  2571 => x"436f6c6f",
  2572 => x"72000000",
  2573 => x"44696666",
  2574 => x"6963756c",
  2575 => x"74792041",
  2576 => x"00000000",
  2577 => x"44696666",
  2578 => x"6963756c",
  2579 => x"74792042",
  2580 => x"00000000",
  2581 => x"53656c65",
  2582 => x"63740000",
  2583 => x"53746172",
  2584 => x"74000000",
  2585 => x"4c6f6164",
  2586 => x"20524f4d",
  2587 => x"20100000",
  2588 => x"45786974",
  2589 => x"00000000",
  2590 => x"524f4d20",
  2591 => x"6c6f6164",
  2592 => x"696e6720",
  2593 => x"6661696c",
  2594 => x"65640000",
  2595 => x"4f4b0000",
  2596 => x"496e6974",
  2597 => x"69616c69",
  2598 => x"7a696e67",
  2599 => x"20534420",
  2600 => x"63617264",
  2601 => x"0a000000",
  2602 => x"16200000",
  2603 => x"14200000",
  2604 => x"15200000",
  2605 => x"53442069",
  2606 => x"6e69742e",
  2607 => x"2e2e0a00",
  2608 => x"53442063",
  2609 => x"61726420",
  2610 => x"72657365",
  2611 => x"74206661",
  2612 => x"696c6564",
  2613 => x"210a0000",
  2614 => x"53444843",
  2615 => x"20657272",
  2616 => x"6f72210a",
  2617 => x"00000000",
  2618 => x"57726974",
  2619 => x"65206661",
  2620 => x"696c6564",
  2621 => x"0a000000",
  2622 => x"52656164",
  2623 => x"20666169",
  2624 => x"6c65640a",
  2625 => x"00000000",
  2626 => x"43617264",
  2627 => x"20696e69",
  2628 => x"74206661",
  2629 => x"696c6564",
  2630 => x"0a000000",
  2631 => x"46415431",
  2632 => x"36202020",
  2633 => x"00000000",
  2634 => x"46415433",
  2635 => x"32202020",
  2636 => x"00000000",
  2637 => x"4e6f2070",
  2638 => x"61727469",
  2639 => x"74696f6e",
  2640 => x"20736967",
  2641 => x"0a000000",
  2642 => x"42616420",
  2643 => x"70617274",
  2644 => x"0a000000",
  2645 => x"4261636b",
  2646 => x"00000000",
  2647 => x"00000002",
  2648 => x"00000002",
  2649 => x"0000280c",
  2650 => x"0000035a",
  2651 => x"00000001",
  2652 => x"00002814",
  2653 => x"00000000",
  2654 => x"00000001",
  2655 => x"00002820",
  2656 => x"00000001",
  2657 => x"00000001",
  2658 => x"0000282c",
  2659 => x"00000002",
  2660 => x"00000001",
  2661 => x"00002834",
  2662 => x"00000003",
  2663 => x"00000001",
  2664 => x"00002844",
  2665 => x"00000004",
  2666 => x"00000002",
  2667 => x"00002854",
  2668 => x"0000036e",
  2669 => x"00000002",
  2670 => x"0000285c",
  2671 => x"00000a3f",
  2672 => x"00000002",
  2673 => x"00002864",
  2674 => x"000027cf",
  2675 => x"00000002",
  2676 => x"00002870",
  2677 => x"000014a6",
  2678 => x"00000000",
  2679 => x"00000000",
  2680 => x"00000000",
  2681 => x"00000004",
  2682 => x"00002878",
  2683 => x"000029e4",
  2684 => x"00000004",
  2685 => x"0000288c",
  2686 => x"00002960",
  2687 => x"00000000",
  2688 => x"00000000",
  2689 => x"00000000",
  2690 => x"00000000",
  2691 => x"00000000",
  2692 => x"00000000",
  2693 => x"00000000",
  2694 => x"00000000",
  2695 => x"00000000",
  2696 => x"00000000",
  2697 => x"00000000",
  2698 => x"00000000",
  2699 => x"00000000",
  2700 => x"00000000",
  2701 => x"00000000",
  2702 => x"00000000",
  2703 => x"00000000",
  2704 => x"00000000",
  2705 => x"00000000",
  2706 => x"00000000",
  2707 => x"00000000",
  2708 => x"00000006",
  2709 => x"00000000",
  2710 => x"00000000",
  2711 => x"00000002",
  2712 => x"00002ec0",
  2713 => x"00002594",
  2714 => x"00000002",
  2715 => x"00002ede",
  2716 => x"00002594",
  2717 => x"00000002",
  2718 => x"00002efc",
  2719 => x"00002594",
  2720 => x"00000002",
  2721 => x"00002f1a",
  2722 => x"00002594",
  2723 => x"00000002",
  2724 => x"00002f38",
  2725 => x"00002594",
  2726 => x"00000002",
  2727 => x"00002f56",
  2728 => x"00002594",
  2729 => x"00000002",
  2730 => x"00002f74",
  2731 => x"00002594",
  2732 => x"00000002",
  2733 => x"00002f92",
  2734 => x"00002594",
  2735 => x"00000002",
  2736 => x"00002fb0",
  2737 => x"00002594",
  2738 => x"00000002",
  2739 => x"00002fce",
  2740 => x"00002594",
  2741 => x"00000002",
  2742 => x"00002fec",
  2743 => x"00002594",
  2744 => x"00000002",
  2745 => x"0000300a",
  2746 => x"00002594",
  2747 => x"00000002",
  2748 => x"00003028",
  2749 => x"00002594",
  2750 => x"00000004",
  2751 => x"00002954",
  2752 => x"00000000",
  2753 => x"00000000",
  2754 => x"00000000",
  2755 => x"00002754",
  2756 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

