-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80e7",
     9 => x"e4080b0b",
    10 => x"80e7e808",
    11 => x"0b0b80e7",
    12 => x"ec080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"e7ec0c0b",
    16 => x"0b80e7e8",
    17 => x"0c0b0b80",
    18 => x"e7e40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80e184",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80e7e470",
    57 => x"80f29827",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51b1bc",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80e7",
    65 => x"f40c9f0b",
    66 => x"80e7f80c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"e7f808ff",
    70 => x"0580e7f8",
    71 => x"0c80e7f8",
    72 => x"088025e8",
    73 => x"3880e7f4",
    74 => x"08ff0580",
    75 => x"e7f40c80",
    76 => x"e7f40880",
    77 => x"25d03880",
    78 => x"0b80e7f8",
    79 => x"0c800b80",
    80 => x"e7f40c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80e7f408",
   100 => x"25913882",
   101 => x"c82d80e7",
   102 => x"f408ff05",
   103 => x"80e7f40c",
   104 => x"838a0480",
   105 => x"e7f40880",
   106 => x"e7f80853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80e7f408",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"e7f80881",
   116 => x"0580e7f8",
   117 => x"0c80e7f8",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80e7f8",
   121 => x"0c80e7f4",
   122 => x"08810580",
   123 => x"e7f40c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480e7",
   128 => x"f8088105",
   129 => x"80e7f80c",
   130 => x"80e7f808",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80e7f8",
   134 => x"0c80e7f4",
   135 => x"08810580",
   136 => x"e7f40c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"e7fc0cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"e7fc0c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280e7",
   177 => x"fc088407",
   178 => x"80e7fc0c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80e4",
   183 => x"840c8171",
   184 => x"2bff05f6",
   185 => x"880cfecc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80e7fc",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80e7",
   208 => x"e40c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"86c72d86",
  1093 => x"c72d86c7",
  1094 => x"2d86c72d",
  1095 => x"86c72d86",
  1096 => x"c72d86c7",
  1097 => x"2d86c72d",
  1098 => x"86c72d86",
  1099 => x"c72d86c7",
  1100 => x"2d86c72d",
  1101 => x"86c72d86",
  1102 => x"c72d86c7",
  1103 => x"2d86c72d",
  1104 => x"86c72d86",
  1105 => x"c72d86c7",
  1106 => x"2d86c72d",
  1107 => x"86c72d86",
  1108 => x"c72d86c7",
  1109 => x"2d86c72d",
  1110 => x"86c72d86",
  1111 => x"c72d86c7",
  1112 => x"2d86c72d",
  1113 => x"86c72d86",
  1114 => x"c72d86c7",
  1115 => x"2d86c72d",
  1116 => x"86c72d86",
  1117 => x"c72d86c7",
  1118 => x"2d86c72d",
  1119 => x"86c72d86",
  1120 => x"c72d86c7",
  1121 => x"2d86c72d",
  1122 => x"86c72d86",
  1123 => x"c72d86c7",
  1124 => x"2d86c72d",
  1125 => x"86c72d86",
  1126 => x"c72d86c7",
  1127 => x"2d86c72d",
  1128 => x"86c72d86",
  1129 => x"c72d86c7",
  1130 => x"2d86c72d",
  1131 => x"86c72d86",
  1132 => x"c72d86c7",
  1133 => x"2d86c72d",
  1134 => x"86c72d86",
  1135 => x"c72d86c7",
  1136 => x"2d86c72d",
  1137 => x"86c72d86",
  1138 => x"c72d86c7",
  1139 => x"2d86c72d",
  1140 => x"86c72d86",
  1141 => x"c72d86c7",
  1142 => x"2d86c72d",
  1143 => x"86c72d86",
  1144 => x"c72d86c7",
  1145 => x"2d86c72d",
  1146 => x"86c72d86",
  1147 => x"c72d86c7",
  1148 => x"2d86c72d",
  1149 => x"86c72d86",
  1150 => x"c72d86c7",
  1151 => x"2d86c72d",
  1152 => x"86c72d86",
  1153 => x"c72d86c7",
  1154 => x"2d86c72d",
  1155 => x"86c72d86",
  1156 => x"c72d86c7",
  1157 => x"2d86c72d",
  1158 => x"86c72d86",
  1159 => x"c72d86c7",
  1160 => x"2d86c72d",
  1161 => x"86c72d86",
  1162 => x"c72d86c7",
  1163 => x"2d86c72d",
  1164 => x"86c72d86",
  1165 => x"c72d86c7",
  1166 => x"2d86c72d",
  1167 => x"86c72d86",
  1168 => x"c72d86c7",
  1169 => x"2d86c72d",
  1170 => x"86c72d86",
  1171 => x"c72d86c7",
  1172 => x"2d86c72d",
  1173 => x"86c72d86",
  1174 => x"c72d86c7",
  1175 => x"2d86c72d",
  1176 => x"86c72d86",
  1177 => x"c72d86c7",
  1178 => x"2d86c72d",
  1179 => x"86c72d86",
  1180 => x"c72d86c7",
  1181 => x"2d86c72d",
  1182 => x"86c72d86",
  1183 => x"c72d86c7",
  1184 => x"2d86c72d",
  1185 => x"86c72d86",
  1186 => x"c72d86c7",
  1187 => x"2d86c72d",
  1188 => x"86c72d86",
  1189 => x"c72d86c7",
  1190 => x"2d86c72d",
  1191 => x"86c72d86",
  1192 => x"c72d86c7",
  1193 => x"2d86c72d",
  1194 => x"86c72d86",
  1195 => x"c72d86c7",
  1196 => x"2d86c72d",
  1197 => x"86c72d86",
  1198 => x"c72d86c7",
  1199 => x"2d86c72d",
  1200 => x"86c72d86",
  1201 => x"c72d86c7",
  1202 => x"2d86c72d",
  1203 => x"86c72d86",
  1204 => x"c72d86c7",
  1205 => x"2d86c72d",
  1206 => x"86c72d86",
  1207 => x"c72d86c7",
  1208 => x"2d86c72d",
  1209 => x"86c72d86",
  1210 => x"c72d86c7",
  1211 => x"2d86c72d",
  1212 => x"86c72d86",
  1213 => x"c72d86c7",
  1214 => x"2d86c72d",
  1215 => x"86c72d86",
  1216 => x"c72d86c7",
  1217 => x"2d86c72d",
  1218 => x"86c72d86",
  1219 => x"c72d86c7",
  1220 => x"2d86c72d",
  1221 => x"86c72d86",
  1222 => x"c72d86c7",
  1223 => x"2d86c72d",
  1224 => x"86c72d86",
  1225 => x"c72d86c7",
  1226 => x"2d86c72d",
  1227 => x"86c72d86",
  1228 => x"c72d86c7",
  1229 => x"2d86c72d",
  1230 => x"86c72d86",
  1231 => x"c72d86c7",
  1232 => x"2d86c72d",
  1233 => x"86c72d86",
  1234 => x"c72d86c7",
  1235 => x"2d86c72d",
  1236 => x"86c72d86",
  1237 => x"c72d86c7",
  1238 => x"2d86c72d",
  1239 => x"86c72d86",
  1240 => x"c72d86c7",
  1241 => x"2d86c72d",
  1242 => x"86c72d86",
  1243 => x"c72d86c7",
  1244 => x"2d86c72d",
  1245 => x"86c72d86",
  1246 => x"c72d86c7",
  1247 => x"2d86c72d",
  1248 => x"86c72d86",
  1249 => x"c72d86c7",
  1250 => x"2d86c72d",
  1251 => x"86c72d86",
  1252 => x"c72d86c7",
  1253 => x"2d86c72d",
  1254 => x"86c72d86",
  1255 => x"c72d86c7",
  1256 => x"2d86c72d",
  1257 => x"86c72d86",
  1258 => x"c72d86c7",
  1259 => x"2d86c72d",
  1260 => x"86c72d86",
  1261 => x"c72d86c7",
  1262 => x"2d86c72d",
  1263 => x"86c72d86",
  1264 => x"c72d86c7",
  1265 => x"2d86c72d",
  1266 => x"86c72d86",
  1267 => x"c72d86c7",
  1268 => x"2d86c72d",
  1269 => x"86c72d86",
  1270 => x"c72d86c7",
  1271 => x"2d86c72d",
  1272 => x"86c72d86",
  1273 => x"c72d86c7",
  1274 => x"2d86c72d",
  1275 => x"86c72d86",
  1276 => x"c72d86c7",
  1277 => x"2d86c72d",
  1278 => x"86c72d86",
  1279 => x"c72d86c7",
  1280 => x"2d86c72d",
  1281 => x"86c72d86",
  1282 => x"c72d86c7",
  1283 => x"2d86c72d",
  1284 => x"86c72d86",
  1285 => x"c72d86c7",
  1286 => x"2d86c72d",
  1287 => x"86c72d86",
  1288 => x"c72d86c7",
  1289 => x"2d86c72d",
  1290 => x"86c72d86",
  1291 => x"c72d86c7",
  1292 => x"2d86c72d",
  1293 => x"86c72d86",
  1294 => x"c72d86c7",
  1295 => x"2d86c72d",
  1296 => x"86c72d86",
  1297 => x"c72d86c7",
  1298 => x"2d86c72d",
  1299 => x"86c72d86",
  1300 => x"c72d86c7",
  1301 => x"2d86c72d",
  1302 => x"86c72d86",
  1303 => x"c72d86c7",
  1304 => x"2d86c72d",
  1305 => x"86c72d86",
  1306 => x"c72d86c7",
  1307 => x"2d86c72d",
  1308 => x"86c72d86",
  1309 => x"c72d86c7",
  1310 => x"2d86c72d",
  1311 => x"86c72d86",
  1312 => x"c72d86c7",
  1313 => x"2d86c72d",
  1314 => x"86c72d86",
  1315 => x"c72d86c7",
  1316 => x"2d86c72d",
  1317 => x"86c72d86",
  1318 => x"c72d86c7",
  1319 => x"2d86c72d",
  1320 => x"86c72d86",
  1321 => x"c72d86c7",
  1322 => x"2d86c72d",
  1323 => x"86c72d86",
  1324 => x"c72d86c7",
  1325 => x"2d86c72d",
  1326 => x"86c72d86",
  1327 => x"c72d86c7",
  1328 => x"2d86c72d",
  1329 => x"86c72d86",
  1330 => x"c72d86c7",
  1331 => x"2d86c72d",
  1332 => x"86c72d86",
  1333 => x"c72d86c7",
  1334 => x"2d86c72d",
  1335 => x"86c72d86",
  1336 => x"c72d86c7",
  1337 => x"2d86c72d",
  1338 => x"86c72d86",
  1339 => x"c72d86c7",
  1340 => x"2d86c72d",
  1341 => x"86c72d86",
  1342 => x"c72d86c7",
  1343 => x"2d86c72d",
  1344 => x"86c72d86",
  1345 => x"c72d86c7",
  1346 => x"2d86c72d",
  1347 => x"86c72d86",
  1348 => x"c72d86c7",
  1349 => x"2d86c72d",
  1350 => x"86c72d86",
  1351 => x"c72d86c7",
  1352 => x"2d86c72d",
  1353 => x"86c72d86",
  1354 => x"c72d86c7",
  1355 => x"2d86c72d",
  1356 => x"86c72d86",
  1357 => x"c72d86c7",
  1358 => x"2d86c72d",
  1359 => x"86c72d86",
  1360 => x"c72d86c7",
  1361 => x"2d86c72d",
  1362 => x"86c72d86",
  1363 => x"c72d86c7",
  1364 => x"2d86c72d",
  1365 => x"86c72d86",
  1366 => x"c72d86c7",
  1367 => x"2d86c72d",
  1368 => x"86c72d86",
  1369 => x"c72d86c7",
  1370 => x"2d86c72d",
  1371 => x"86c72d86",
  1372 => x"c72d86c7",
  1373 => x"2d86c72d",
  1374 => x"86c72d86",
  1375 => x"c72d86c7",
  1376 => x"2d86c72d",
  1377 => x"86c72d86",
  1378 => x"c72d86c7",
  1379 => x"2d86c72d",
  1380 => x"86c72d86",
  1381 => x"c72d86c7",
  1382 => x"2d86c72d",
  1383 => x"86c72d86",
  1384 => x"c72d86c7",
  1385 => x"2d86c72d",
  1386 => x"86c72d86",
  1387 => x"c72d86c7",
  1388 => x"2d86c72d",
  1389 => x"86c72d86",
  1390 => x"c72d86c7",
  1391 => x"2d86c72d",
  1392 => x"86c72d86",
  1393 => x"c72d86c7",
  1394 => x"2d86c72d",
  1395 => x"86c72d86",
  1396 => x"c72d86c7",
  1397 => x"2d86c72d",
  1398 => x"86c72d86",
  1399 => x"c72d86c7",
  1400 => x"2d86c72d",
  1401 => x"86c72d86",
  1402 => x"c72d86c7",
  1403 => x"2d86c72d",
  1404 => x"86c72d86",
  1405 => x"c72d86c7",
  1406 => x"2d86c72d",
  1407 => x"86c72d86",
  1408 => x"c72d86c7",
  1409 => x"2d86c72d",
  1410 => x"86c72d86",
  1411 => x"c72d86c7",
  1412 => x"2d86c72d",
  1413 => x"86c72d86",
  1414 => x"c72d86c7",
  1415 => x"2d86c72d",
  1416 => x"86c72d86",
  1417 => x"c72d86c7",
  1418 => x"2d86c72d",
  1419 => x"86c72d86",
  1420 => x"c72d86c7",
  1421 => x"2d86c72d",
  1422 => x"86c72d86",
  1423 => x"c72d86c7",
  1424 => x"2d86c72d",
  1425 => x"86c72d86",
  1426 => x"c72d86c7",
  1427 => x"2d86c72d",
  1428 => x"86c72d86",
  1429 => x"c72d86c7",
  1430 => x"2d86c72d",
  1431 => x"86c72d86",
  1432 => x"c72d86c7",
  1433 => x"2d86c72d",
  1434 => x"86c72d86",
  1435 => x"c72d86c7",
  1436 => x"2d86c72d",
  1437 => x"86c72d86",
  1438 => x"c72d86c7",
  1439 => x"2d86c72d",
  1440 => x"86c72d86",
  1441 => x"c72d86c7",
  1442 => x"2d86c72d",
  1443 => x"86c72d86",
  1444 => x"c72d86c7",
  1445 => x"2d86c72d",
  1446 => x"86c72d86",
  1447 => x"c72d86c7",
  1448 => x"2d86c72d",
  1449 => x"86c72d86",
  1450 => x"c72d86c7",
  1451 => x"2d86c72d",
  1452 => x"86c72d86",
  1453 => x"c72d86c7",
  1454 => x"2d86c72d",
  1455 => x"86c72d86",
  1456 => x"c72d86c7",
  1457 => x"2d86c72d",
  1458 => x"86c72d86",
  1459 => x"c72d86c7",
  1460 => x"2d86c72d",
  1461 => x"86c72d86",
  1462 => x"c72d86c7",
  1463 => x"2d86c72d",
  1464 => x"86c72d86",
  1465 => x"c72d86c7",
  1466 => x"2d86c72d",
  1467 => x"86c72d86",
  1468 => x"c72d86c7",
  1469 => x"2d86c72d",
  1470 => x"86c72d86",
  1471 => x"c72d86c7",
  1472 => x"2d86c72d",
  1473 => x"86c72d86",
  1474 => x"c72d86c7",
  1475 => x"2d86c72d",
  1476 => x"86c72d86",
  1477 => x"c72d86c7",
  1478 => x"2d86c72d",
  1479 => x"86c72d86",
  1480 => x"c72d86c7",
  1481 => x"2d86c72d",
  1482 => x"86c72d86",
  1483 => x"c72d86c7",
  1484 => x"2d86c72d",
  1485 => x"86c72d86",
  1486 => x"c72d86c7",
  1487 => x"2d86c72d",
  1488 => x"86c72d86",
  1489 => x"c72d86c7",
  1490 => x"2d86c72d",
  1491 => x"86c72d86",
  1492 => x"c72d86c7",
  1493 => x"2d86c72d",
  1494 => x"86c72d86",
  1495 => x"c72d86c7",
  1496 => x"2d86c72d",
  1497 => x"86c72d86",
  1498 => x"c72d86c7",
  1499 => x"2d86c72d",
  1500 => x"86c72d86",
  1501 => x"c72d86c7",
  1502 => x"2d86c72d",
  1503 => x"86c72d86",
  1504 => x"c72d86c7",
  1505 => x"2d86c72d",
  1506 => x"86c72d86",
  1507 => x"c72d86c7",
  1508 => x"2d86c72d",
  1509 => x"86c72d86",
  1510 => x"c72d86c7",
  1511 => x"2d86c72d",
  1512 => x"86c72d86",
  1513 => x"c72d86c7",
  1514 => x"2d86c72d",
  1515 => x"86c72d86",
  1516 => x"c72d86c7",
  1517 => x"2d86c72d",
  1518 => x"86c72d86",
  1519 => x"c72d86c7",
  1520 => x"2d86c72d",
  1521 => x"86c72d86",
  1522 => x"c72d86c7",
  1523 => x"2d86c72d",
  1524 => x"0402dc05",
  1525 => x"0d7a5380",
  1526 => x"59810bec",
  1527 => x"0c840bec",
  1528 => x"0c725280",
  1529 => x"e8805180",
  1530 => x"d7ce2d80",
  1531 => x"e7e40879",
  1532 => x"2e819f38",
  1533 => x"80e88408",
  1534 => x"79ff1256",
  1535 => x"59557485",
  1536 => x"2e098106",
  1537 => x"a4387251",
  1538 => x"86a02da2",
  1539 => x"902da290",
  1540 => x"2da2902d",
  1541 => x"a2902da2",
  1542 => x"902da290",
  1543 => x"2d80e488",
  1544 => x"51bafa2d",
  1545 => x"8153b1b2",
  1546 => x"0473802e",
  1547 => x"8b388118",
  1548 => x"74812a55",
  1549 => x"58b0a904",
  1550 => x"f7185881",
  1551 => x"59807525",
  1552 => x"80d03877",
  1553 => x"52735184",
  1554 => x"a82d80e8",
  1555 => x"d05280e8",
  1556 => x"805180da",
  1557 => x"a42d80e7",
  1558 => x"e408802e",
  1559 => x"9b3880e8",
  1560 => x"d05783fc",
  1561 => x"56767084",
  1562 => x"055808e8",
  1563 => x"0cfc1656",
  1564 => x"758025f1",
  1565 => x"38b18004",
  1566 => x"80e7e408",
  1567 => x"59848055",
  1568 => x"80e88051",
  1569 => x"80d9f32d",
  1570 => x"fc801581",
  1571 => x"155555b0",
  1572 => x"bd0480e8",
  1573 => x"8408f80c",
  1574 => x"805186da",
  1575 => x"2d78802e",
  1576 => x"883880e4",
  1577 => x"8851b1ad",
  1578 => x"0480e58c",
  1579 => x"51bafa2d",
  1580 => x"78537280",
  1581 => x"e7e40c02",
  1582 => x"a4050d04",
  1583 => x"02ec050d",
  1584 => x"840bec0c",
  1585 => x"b8a92db4",
  1586 => x"de2d81f9",
  1587 => x"2d8353b8",
  1588 => x"8c2d8151",
  1589 => x"858d2dff",
  1590 => x"13537280",
  1591 => x"25f13884",
  1592 => x"0bec0c80",
  1593 => x"e2b85186",
  1594 => x"a02d80cd",
  1595 => x"ee2d80e7",
  1596 => x"e408802e",
  1597 => x"82d13881",
  1598 => x"0bec0c84",
  1599 => x"0bec0c80",
  1600 => x"e1945280",
  1601 => x"e8805180",
  1602 => x"d7ce2d80",
  1603 => x"e7e40880",
  1604 => x"2e80cc38",
  1605 => x"80e8d052",
  1606 => x"80e88051",
  1607 => x"80daa42d",
  1608 => x"80e7e408",
  1609 => x"802eb838",
  1610 => x"80e8d00b",
  1611 => x"80f52d80",
  1612 => x"e6900c80",
  1613 => x"e8d10b80",
  1614 => x"f52d80e6",
  1615 => x"940c80e8",
  1616 => x"d20b80f5",
  1617 => x"2d80e698",
  1618 => x"0c80e8d3",
  1619 => x"0b80f52d",
  1620 => x"80e69c0c",
  1621 => x"80e8d40b",
  1622 => x"80f52d80",
  1623 => x"e6a00c80",
  1624 => x"e1a45280",
  1625 => x"e8805180",
  1626 => x"d7ce2d80",
  1627 => x"e7e40880",
  1628 => x"2e80cc38",
  1629 => x"80e8d052",
  1630 => x"80e88051",
  1631 => x"80daa42d",
  1632 => x"80e7e408",
  1633 => x"802eb838",
  1634 => x"80e8d00b",
  1635 => x"80f52d80",
  1636 => x"e5fc0c80",
  1637 => x"e8d10b80",
  1638 => x"f52d80e6",
  1639 => x"800c80e8",
  1640 => x"d20b80f5",
  1641 => x"2d80e684",
  1642 => x"0c80e8d3",
  1643 => x"0b80f52d",
  1644 => x"80e6880c",
  1645 => x"80e8d40b",
  1646 => x"80f52d80",
  1647 => x"e68c0caf",
  1648 => x"d15180e0",
  1649 => x"fb2d80e4",
  1650 => x"8851bafa",
  1651 => x"2db8cb2d",
  1652 => x"b4ea2dbb",
  1653 => x"8d2d80e4",
  1654 => x"9c0b80f5",
  1655 => x"2d80e5f8",
  1656 => x"08708106",
  1657 => x"55565472",
  1658 => x"802e8538",
  1659 => x"73840754",
  1660 => x"74812a70",
  1661 => x"81065153",
  1662 => x"72802e85",
  1663 => x"38738207",
  1664 => x"5474822a",
  1665 => x"70810651",
  1666 => x"5372802e",
  1667 => x"85387381",
  1668 => x"07547483",
  1669 => x"2a708106",
  1670 => x"51537280",
  1671 => x"2e853873",
  1672 => x"88075474",
  1673 => x"842a7081",
  1674 => x"06515372",
  1675 => x"802e8538",
  1676 => x"73900754",
  1677 => x"73fc0c86",
  1678 => x"5380e7e4",
  1679 => x"08833884",
  1680 => x"5372ec0c",
  1681 => x"b3d00480",
  1682 => x"0b80e7e4",
  1683 => x"0c029405",
  1684 => x"0d047198",
  1685 => x"0c04ffb0",
  1686 => x"0880e7e4",
  1687 => x"0c04810b",
  1688 => x"ffb00c04",
  1689 => x"800bffb0",
  1690 => x"0c0402f4",
  1691 => x"050db5f8",
  1692 => x"0480e7e4",
  1693 => x"0881f02e",
  1694 => x"0981068a",
  1695 => x"38810b80",
  1696 => x"e5f00cb5",
  1697 => x"f80480e7",
  1698 => x"e40881e0",
  1699 => x"2e098106",
  1700 => x"8a38810b",
  1701 => x"80e5f40c",
  1702 => x"b5f80480",
  1703 => x"e7e40852",
  1704 => x"80e5f408",
  1705 => x"802e8938",
  1706 => x"80e7e408",
  1707 => x"81800552",
  1708 => x"71842c72",
  1709 => x"8f065353",
  1710 => x"80e5f008",
  1711 => x"802e9a38",
  1712 => x"72842980",
  1713 => x"e5b00572",
  1714 => x"1381712b",
  1715 => x"70097308",
  1716 => x"06730c51",
  1717 => x"5353b5ec",
  1718 => x"04728429",
  1719 => x"80e5b005",
  1720 => x"72138371",
  1721 => x"2b720807",
  1722 => x"720c5353",
  1723 => x"800b80e5",
  1724 => x"f40c800b",
  1725 => x"80e5f00c",
  1726 => x"80e88c51",
  1727 => x"b6ff2d80",
  1728 => x"e7e408ff",
  1729 => x"24feea38",
  1730 => x"800b80e7",
  1731 => x"e40c028c",
  1732 => x"050d0402",
  1733 => x"f8050d80",
  1734 => x"e5b0528f",
  1735 => x"51807270",
  1736 => x"8405540c",
  1737 => x"ff115170",
  1738 => x"8025f238",
  1739 => x"0288050d",
  1740 => x"0402f005",
  1741 => x"0d7551b4",
  1742 => x"e42d7082",
  1743 => x"2cfc0680",
  1744 => x"e5b01172",
  1745 => x"109e0671",
  1746 => x"0870722a",
  1747 => x"70830682",
  1748 => x"742b7009",
  1749 => x"7406760c",
  1750 => x"54515657",
  1751 => x"535153b4",
  1752 => x"de2d7180",
  1753 => x"e7e40c02",
  1754 => x"90050d04",
  1755 => x"02fc050d",
  1756 => x"72518071",
  1757 => x"0c800b84",
  1758 => x"120c0284",
  1759 => x"050d0402",
  1760 => x"f0050d75",
  1761 => x"70088412",
  1762 => x"08535353",
  1763 => x"ff547171",
  1764 => x"2ea838b4",
  1765 => x"e42d8413",
  1766 => x"08708429",
  1767 => x"14881170",
  1768 => x"087081ff",
  1769 => x"06841808",
  1770 => x"81118706",
  1771 => x"841a0c53",
  1772 => x"51555151",
  1773 => x"51b4de2d",
  1774 => x"71547380",
  1775 => x"e7e40c02",
  1776 => x"90050d04",
  1777 => x"02f8050d",
  1778 => x"b4e42de0",
  1779 => x"08708b2a",
  1780 => x"70810651",
  1781 => x"52527080",
  1782 => x"2ea13880",
  1783 => x"e88c0870",
  1784 => x"842980e8",
  1785 => x"94057381",
  1786 => x"ff06710c",
  1787 => x"515180e8",
  1788 => x"8c088111",
  1789 => x"870680e8",
  1790 => x"8c0c5180",
  1791 => x"0b80e8b4",
  1792 => x"0cb4d62d",
  1793 => x"b4de2d02",
  1794 => x"88050d04",
  1795 => x"02fc050d",
  1796 => x"b4e42d81",
  1797 => x"0b80e8b4",
  1798 => x"0cb4de2d",
  1799 => x"80e8b408",
  1800 => x"5170f938",
  1801 => x"0284050d",
  1802 => x"0402fc05",
  1803 => x"0d80e88c",
  1804 => x"51b6ec2d",
  1805 => x"b6932db7",
  1806 => x"c451b4d2",
  1807 => x"2d028405",
  1808 => x"0d0480e8",
  1809 => x"bc0880e7",
  1810 => x"e40c0402",
  1811 => x"fc050d81",
  1812 => x"0b80e6a4",
  1813 => x"0c815185",
  1814 => x"8d2d0284",
  1815 => x"050d0402",
  1816 => x"fc050db8",
  1817 => x"e904b4ea",
  1818 => x"2d80f651",
  1819 => x"b6b12d80",
  1820 => x"e7e408f2",
  1821 => x"3880da51",
  1822 => x"b6b12d80",
  1823 => x"e7e408e6",
  1824 => x"3880e6a0",
  1825 => x"0851b6b1",
  1826 => x"2d80e7e4",
  1827 => x"08d83880",
  1828 => x"e7e40880",
  1829 => x"e6a40c80",
  1830 => x"e7e40851",
  1831 => x"858d2d02",
  1832 => x"84050d04",
  1833 => x"02ec050d",
  1834 => x"76548052",
  1835 => x"870b8815",
  1836 => x"80f52d56",
  1837 => x"53747224",
  1838 => x"8338a053",
  1839 => x"72518384",
  1840 => x"2d81128b",
  1841 => x"1580f52d",
  1842 => x"54527272",
  1843 => x"25de3802",
  1844 => x"94050d04",
  1845 => x"02f0050d",
  1846 => x"80e8bc08",
  1847 => x"5481f92d",
  1848 => x"800b80e8",
  1849 => x"c00c7308",
  1850 => x"802e8189",
  1851 => x"38820b80",
  1852 => x"e7f80c80",
  1853 => x"e8c0088f",
  1854 => x"0680e7f4",
  1855 => x"0c730852",
  1856 => x"71832e96",
  1857 => x"38718326",
  1858 => x"89387181",
  1859 => x"2eb038ba",
  1860 => x"de047185",
  1861 => x"2ea038ba",
  1862 => x"de048814",
  1863 => x"80f52d84",
  1864 => x"150880e2",
  1865 => x"d0535452",
  1866 => x"86a02d71",
  1867 => x"84291370",
  1868 => x"085252ba",
  1869 => x"e2047351",
  1870 => x"b9a42dba",
  1871 => x"de0480e5",
  1872 => x"f8088815",
  1873 => x"082c7081",
  1874 => x"06515271",
  1875 => x"802e8838",
  1876 => x"80e2d451",
  1877 => x"badb0480",
  1878 => x"e2d85186",
  1879 => x"a02d8414",
  1880 => x"085186a0",
  1881 => x"2d80e8c0",
  1882 => x"08810580",
  1883 => x"e8c00c8c",
  1884 => x"1454b9e6",
  1885 => x"04029005",
  1886 => x"0d047180",
  1887 => x"e8bc0cb9",
  1888 => x"d42d80e8",
  1889 => x"c008ff05",
  1890 => x"80e8c40c",
  1891 => x"0402e805",
  1892 => x"0d80e8bc",
  1893 => x"0880e8c8",
  1894 => x"08575580",
  1895 => x"f651b6b1",
  1896 => x"2d80e7e4",
  1897 => x"08812a70",
  1898 => x"81065152",
  1899 => x"71802ea2",
  1900 => x"38bbb704",
  1901 => x"b4ea2d80",
  1902 => x"f651b6b1",
  1903 => x"2d80e7e4",
  1904 => x"08f23880",
  1905 => x"e6a40881",
  1906 => x"327080e6",
  1907 => x"a40c5185",
  1908 => x"8d2d800b",
  1909 => x"80e8b80c",
  1910 => x"8c51b6b1",
  1911 => x"2d80e7e4",
  1912 => x"08812a70",
  1913 => x"81065152",
  1914 => x"71802e80",
  1915 => x"d33880e5",
  1916 => x"fc0880e6",
  1917 => x"900880e5",
  1918 => x"fc0c80e6",
  1919 => x"900c80e6",
  1920 => x"800880e6",
  1921 => x"940880e6",
  1922 => x"800c80e6",
  1923 => x"940c80e6",
  1924 => x"840880e6",
  1925 => x"980880e6",
  1926 => x"840c80e6",
  1927 => x"980c80e6",
  1928 => x"880880e6",
  1929 => x"9c0880e6",
  1930 => x"880c80e6",
  1931 => x"9c0c80e6",
  1932 => x"8c0880e6",
  1933 => x"a00880e6",
  1934 => x"8c0c7080",
  1935 => x"e6a00c52",
  1936 => x"80e6a408",
  1937 => x"82943880",
  1938 => x"e6900851",
  1939 => x"b6b12d80",
  1940 => x"e7e40880",
  1941 => x"2e8b3880",
  1942 => x"e8b80881",
  1943 => x"0780e8b8",
  1944 => x"0c80e694",
  1945 => x"0851b6b1",
  1946 => x"2d80e7e4",
  1947 => x"08802e8b",
  1948 => x"3880e8b8",
  1949 => x"08820780",
  1950 => x"e8b80c80",
  1951 => x"e6980851",
  1952 => x"b6b12d80",
  1953 => x"e7e40880",
  1954 => x"2e8b3880",
  1955 => x"e8b80884",
  1956 => x"0780e8b8",
  1957 => x"0c80e69c",
  1958 => x"0851b6b1",
  1959 => x"2d80e7e4",
  1960 => x"08802e8b",
  1961 => x"3880e8b8",
  1962 => x"08880780",
  1963 => x"e8b80c80",
  1964 => x"e6a00851",
  1965 => x"b6b12d80",
  1966 => x"e7e40880",
  1967 => x"2e8b3880",
  1968 => x"e8b80890",
  1969 => x"0780e8b8",
  1970 => x"0c80e5fc",
  1971 => x"0851b6b1",
  1972 => x"2d80e7e4",
  1973 => x"08802e8c",
  1974 => x"3880e8b8",
  1975 => x"08828007",
  1976 => x"80e8b80c",
  1977 => x"80e68008",
  1978 => x"51b6b12d",
  1979 => x"80e7e408",
  1980 => x"802e8c38",
  1981 => x"80e8b808",
  1982 => x"84800780",
  1983 => x"e8b80c80",
  1984 => x"e6840851",
  1985 => x"b6b12d80",
  1986 => x"e7e40880",
  1987 => x"2e8c3880",
  1988 => x"e8b80888",
  1989 => x"800780e8",
  1990 => x"b80c80e6",
  1991 => x"880851b6",
  1992 => x"b12d80e7",
  1993 => x"e408802e",
  1994 => x"8c3880e8",
  1995 => x"b8089080",
  1996 => x"0780e8b8",
  1997 => x"0c80e68c",
  1998 => x"0851b6b1",
  1999 => x"2d80e7e4",
  2000 => x"08802e8c",
  2001 => x"3880e8b8",
  2002 => x"08a08007",
  2003 => x"80e8b80c",
  2004 => x"80e8b808",
  2005 => x"ed0c80c5",
  2006 => x"a70481f5",
  2007 => x"51b6b12d",
  2008 => x"80e7e408",
  2009 => x"812a7081",
  2010 => x"06515271",
  2011 => x"993880e6",
  2012 => x"900851b6",
  2013 => x"b12d80e7",
  2014 => x"e408812a",
  2015 => x"70810651",
  2016 => x"5271802e",
  2017 => x"b33880e8",
  2018 => x"c4085271",
  2019 => x"802e8a38",
  2020 => x"ff1280e8",
  2021 => x"c40cbfb8",
  2022 => x"0480e8c0",
  2023 => x"081080e8",
  2024 => x"c0080570",
  2025 => x"84291651",
  2026 => x"52881208",
  2027 => x"802e8938",
  2028 => x"ff518812",
  2029 => x"0852712d",
  2030 => x"81f251b6",
  2031 => x"b12d80e7",
  2032 => x"e408812a",
  2033 => x"70810651",
  2034 => x"52719938",
  2035 => x"80e69408",
  2036 => x"51b6b12d",
  2037 => x"80e7e408",
  2038 => x"812a7081",
  2039 => x"06515271",
  2040 => x"802eb538",
  2041 => x"80e8c008",
  2042 => x"ff1180e8",
  2043 => x"c4085653",
  2044 => x"53737225",
  2045 => x"8b388114",
  2046 => x"80e8c40c",
  2047 => x"80c09804",
  2048 => x"72101370",
  2049 => x"84291651",
  2050 => x"52881208",
  2051 => x"802e8938",
  2052 => x"fe518812",
  2053 => x"0852712d",
  2054 => x"81fd51b6",
  2055 => x"b12d80e7",
  2056 => x"e408812a",
  2057 => x"70810651",
  2058 => x"52719938",
  2059 => x"80e69808",
  2060 => x"51b6b12d",
  2061 => x"80e7e408",
  2062 => x"812a7081",
  2063 => x"06515271",
  2064 => x"802eb238",
  2065 => x"80e8c408",
  2066 => x"802e8b38",
  2067 => x"800b80e8",
  2068 => x"c40c80c0",
  2069 => x"f50480e8",
  2070 => x"c0081080",
  2071 => x"e8c00805",
  2072 => x"70842916",
  2073 => x"51528812",
  2074 => x"08802e89",
  2075 => x"38fd5188",
  2076 => x"12085271",
  2077 => x"2d81fa51",
  2078 => x"b6b12d80",
  2079 => x"e7e40881",
  2080 => x"2a708106",
  2081 => x"51527199",
  2082 => x"3880e69c",
  2083 => x"0851b6b1",
  2084 => x"2d80e7e4",
  2085 => x"08812a70",
  2086 => x"81065152",
  2087 => x"71802eb2",
  2088 => x"3880e8c0",
  2089 => x"08ff1154",
  2090 => x"5280e8c4",
  2091 => x"0873258a",
  2092 => x"387280e8",
  2093 => x"c40c80c1",
  2094 => x"d2047110",
  2095 => x"12708429",
  2096 => x"16515288",
  2097 => x"1208802e",
  2098 => x"8938fc51",
  2099 => x"88120852",
  2100 => x"712d80e8",
  2101 => x"c4087053",
  2102 => x"5473802e",
  2103 => x"8b388c15",
  2104 => x"ff155555",
  2105 => x"80c1d904",
  2106 => x"820b80e7",
  2107 => x"f80c718f",
  2108 => x"0680e7f4",
  2109 => x"0c81eb51",
  2110 => x"b6b12d80",
  2111 => x"e7e40881",
  2112 => x"2a708106",
  2113 => x"51527180",
  2114 => x"2ead3874",
  2115 => x"08852e09",
  2116 => x"8106a438",
  2117 => x"881580f5",
  2118 => x"2dff0552",
  2119 => x"71881681",
  2120 => x"b72d7198",
  2121 => x"2b527180",
  2122 => x"25883880",
  2123 => x"0b881681",
  2124 => x"b72d7451",
  2125 => x"b9a42d81",
  2126 => x"f451b6b1",
  2127 => x"2d80e7e4",
  2128 => x"08812a70",
  2129 => x"81065152",
  2130 => x"71802eb3",
  2131 => x"38740885",
  2132 => x"2e098106",
  2133 => x"aa388815",
  2134 => x"80f52d81",
  2135 => x"05527188",
  2136 => x"1681b72d",
  2137 => x"7181ff06",
  2138 => x"8b1680f5",
  2139 => x"2d545272",
  2140 => x"72278738",
  2141 => x"72881681",
  2142 => x"b72d7451",
  2143 => x"b9a42d80",
  2144 => x"da51b6b1",
  2145 => x"2d80e7e4",
  2146 => x"08812a70",
  2147 => x"81065152",
  2148 => x"719a3880",
  2149 => x"e6a00851",
  2150 => x"b6b12d80",
  2151 => x"e7e40881",
  2152 => x"2a708106",
  2153 => x"51527180",
  2154 => x"2e81b338",
  2155 => x"80e8bc08",
  2156 => x"80e8c408",
  2157 => x"55537380",
  2158 => x"2e8b388c",
  2159 => x"13ff1555",
  2160 => x"5380c3b6",
  2161 => x"04720852",
  2162 => x"71822ea8",
  2163 => x"38718226",
  2164 => x"8a387181",
  2165 => x"2ead3880",
  2166 => x"c4de0471",
  2167 => x"832eb738",
  2168 => x"71842e09",
  2169 => x"810680f6",
  2170 => x"38881308",
  2171 => x"51bafa2d",
  2172 => x"80c4de04",
  2173 => x"80e8c408",
  2174 => x"51881308",
  2175 => x"52712d80",
  2176 => x"c4de0481",
  2177 => x"0b881408",
  2178 => x"2b80e5f8",
  2179 => x"083280e5",
  2180 => x"f80c80c4",
  2181 => x"b1048813",
  2182 => x"80f52d81",
  2183 => x"058b1480",
  2184 => x"f52d5354",
  2185 => x"71742483",
  2186 => x"38805473",
  2187 => x"881481b7",
  2188 => x"2db9d42d",
  2189 => x"80c4de04",
  2190 => x"7508802e",
  2191 => x"a4387508",
  2192 => x"51b6b12d",
  2193 => x"80e7e408",
  2194 => x"81065271",
  2195 => x"802e8c38",
  2196 => x"80e8c408",
  2197 => x"51841608",
  2198 => x"52712d88",
  2199 => x"165675d8",
  2200 => x"38805480",
  2201 => x"0b80e7f8",
  2202 => x"0c738f06",
  2203 => x"80e7f40c",
  2204 => x"a0527380",
  2205 => x"e8c4082e",
  2206 => x"09810699",
  2207 => x"3880e8c0",
  2208 => x"08ff0574",
  2209 => x"32700981",
  2210 => x"05707207",
  2211 => x"9f2a9171",
  2212 => x"31515153",
  2213 => x"53715183",
  2214 => x"842d8114",
  2215 => x"548e7425",
  2216 => x"c23880e6",
  2217 => x"a4085271",
  2218 => x"80e7e40c",
  2219 => x"0298050d",
  2220 => x"0402f405",
  2221 => x"0dd45281",
  2222 => x"ff720c71",
  2223 => x"085381ff",
  2224 => x"720c7288",
  2225 => x"2b83fe80",
  2226 => x"06720870",
  2227 => x"81ff0651",
  2228 => x"525381ff",
  2229 => x"720c7271",
  2230 => x"07882b72",
  2231 => x"087081ff",
  2232 => x"06515253",
  2233 => x"81ff720c",
  2234 => x"72710788",
  2235 => x"2b720870",
  2236 => x"81ff0672",
  2237 => x"0780e7e4",
  2238 => x"0c525302",
  2239 => x"8c050d04",
  2240 => x"02f4050d",
  2241 => x"74767181",
  2242 => x"ff06d40c",
  2243 => x"535380e8",
  2244 => x"cc088538",
  2245 => x"71892b52",
  2246 => x"71982ad4",
  2247 => x"0c71902a",
  2248 => x"7081ff06",
  2249 => x"d40c5171",
  2250 => x"882a7081",
  2251 => x"ff06d40c",
  2252 => x"517181ff",
  2253 => x"06d40c72",
  2254 => x"902a7081",
  2255 => x"ff06d40c",
  2256 => x"51d40870",
  2257 => x"81ff0651",
  2258 => x"5182b8bf",
  2259 => x"527081ff",
  2260 => x"2e098106",
  2261 => x"943881ff",
  2262 => x"0bd40cd4",
  2263 => x"087081ff",
  2264 => x"06ff1454",
  2265 => x"515171e5",
  2266 => x"387080e7",
  2267 => x"e40c028c",
  2268 => x"050d0402",
  2269 => x"fc050d81",
  2270 => x"c75181ff",
  2271 => x"0bd40cff",
  2272 => x"11517080",
  2273 => x"25f43802",
  2274 => x"84050d04",
  2275 => x"02f4050d",
  2276 => x"81ff0bd4",
  2277 => x"0c935380",
  2278 => x"5287fc80",
  2279 => x"c15180c6",
  2280 => x"802d80e7",
  2281 => x"e4088c38",
  2282 => x"81ff0bd4",
  2283 => x"0c815380",
  2284 => x"c7bd0480",
  2285 => x"c6f32dff",
  2286 => x"135372db",
  2287 => x"387280e7",
  2288 => x"e40c028c",
  2289 => x"050d0402",
  2290 => x"ec050d81",
  2291 => x"0b80e8cc",
  2292 => x"0c8454d0",
  2293 => x"08708f2a",
  2294 => x"70810651",
  2295 => x"515372f3",
  2296 => x"3872d00c",
  2297 => x"80c6f32d",
  2298 => x"80e2dc51",
  2299 => x"86a02dd0",
  2300 => x"08708f2a",
  2301 => x"70810651",
  2302 => x"515372f3",
  2303 => x"38810bd0",
  2304 => x"0cb15380",
  2305 => x"5284d480",
  2306 => x"c05180c6",
  2307 => x"802d80e7",
  2308 => x"e408812e",
  2309 => x"94387282",
  2310 => x"2e80c438",
  2311 => x"ff135372",
  2312 => x"e238ff14",
  2313 => x"5473ffab",
  2314 => x"3880c6f3",
  2315 => x"2d83aa52",
  2316 => x"849c80c8",
  2317 => x"5180c680",
  2318 => x"2d80e7e4",
  2319 => x"08812e09",
  2320 => x"81069438",
  2321 => x"80c5b12d",
  2322 => x"80e7e408",
  2323 => x"83ffff06",
  2324 => x"537283aa",
  2325 => x"2ea33880",
  2326 => x"c78c2d80",
  2327 => x"c8f30480",
  2328 => x"e2e85186",
  2329 => x"a02d8053",
  2330 => x"80cad104",
  2331 => x"80e38051",
  2332 => x"86a02d80",
  2333 => x"5480caa1",
  2334 => x"0481ff0b",
  2335 => x"d40cb154",
  2336 => x"80c6f32d",
  2337 => x"8fcf5380",
  2338 => x"5287fc80",
  2339 => x"f75180c6",
  2340 => x"802d80e7",
  2341 => x"e4085580",
  2342 => x"e7e40881",
  2343 => x"2e098106",
  2344 => x"9e3881ff",
  2345 => x"0bd40c82",
  2346 => x"0a52849c",
  2347 => x"80e95180",
  2348 => x"c6802d80",
  2349 => x"e7e40880",
  2350 => x"2e8f3880",
  2351 => x"c6f32dff",
  2352 => x"135372c3",
  2353 => x"3880ca94",
  2354 => x"0481ff0b",
  2355 => x"d40c80e7",
  2356 => x"e4085287",
  2357 => x"fc80fa51",
  2358 => x"80c6802d",
  2359 => x"80e7e408",
  2360 => x"b33881ff",
  2361 => x"0bd40cd4",
  2362 => x"085381ff",
  2363 => x"0bd40c81",
  2364 => x"ff0bd40c",
  2365 => x"81ff0bd4",
  2366 => x"0c81ff0b",
  2367 => x"d40c7286",
  2368 => x"2a708106",
  2369 => x"76565153",
  2370 => x"72973880",
  2371 => x"e7e40854",
  2372 => x"80caa104",
  2373 => x"73822efe",
  2374 => x"d338ff14",
  2375 => x"5473fee0",
  2376 => x"387380e8",
  2377 => x"cc0c738c",
  2378 => x"38815287",
  2379 => x"fc80d051",
  2380 => x"80c6802d",
  2381 => x"81ff0bd4",
  2382 => x"0cd00870",
  2383 => x"8f2a7081",
  2384 => x"06515153",
  2385 => x"72f33872",
  2386 => x"d00c81ff",
  2387 => x"0bd40c81",
  2388 => x"537280e7",
  2389 => x"e40c0294",
  2390 => x"050d0402",
  2391 => x"e8050d78",
  2392 => x"55805681",
  2393 => x"ff0bd40c",
  2394 => x"d008708f",
  2395 => x"2a708106",
  2396 => x"51515372",
  2397 => x"f3388281",
  2398 => x"0bd00c81",
  2399 => x"ff0bd40c",
  2400 => x"775287fc",
  2401 => x"80d15180",
  2402 => x"c6802d80",
  2403 => x"dbc6df54",
  2404 => x"80e7e408",
  2405 => x"802e8c38",
  2406 => x"80e3a051",
  2407 => x"86a02d80",
  2408 => x"cbf90481",
  2409 => x"ff0bd40c",
  2410 => x"d4087081",
  2411 => x"ff065153",
  2412 => x"7281fe2e",
  2413 => x"098106a0",
  2414 => x"3880ff53",
  2415 => x"80c5b12d",
  2416 => x"80e7e408",
  2417 => x"75708405",
  2418 => x"570cff13",
  2419 => x"53728025",
  2420 => x"eb388156",
  2421 => x"80cbde04",
  2422 => x"ff145473",
  2423 => x"c63881ff",
  2424 => x"0bd40c81",
  2425 => x"ff0bd40c",
  2426 => x"d008708f",
  2427 => x"2a708106",
  2428 => x"51515372",
  2429 => x"f33872d0",
  2430 => x"0c7580e7",
  2431 => x"e40c0298",
  2432 => x"050d0402",
  2433 => x"e8050d77",
  2434 => x"797b5855",
  2435 => x"55805372",
  2436 => x"7625a538",
  2437 => x"74708105",
  2438 => x"5680f52d",
  2439 => x"74708105",
  2440 => x"5680f52d",
  2441 => x"52527171",
  2442 => x"2e873881",
  2443 => x"5180ccba",
  2444 => x"04811353",
  2445 => x"80cc8f04",
  2446 => x"80517080",
  2447 => x"e7e40c02",
  2448 => x"98050d04",
  2449 => x"02ec050d",
  2450 => x"76557480",
  2451 => x"2e80c438",
  2452 => x"9a1580e0",
  2453 => x"2d5180da",
  2454 => x"ff2d80e7",
  2455 => x"e40880e7",
  2456 => x"e40880ef",
  2457 => x"800c80e7",
  2458 => x"e4085454",
  2459 => x"80eedc08",
  2460 => x"802e9b38",
  2461 => x"941580e0",
  2462 => x"2d5180da",
  2463 => x"ff2d80e7",
  2464 => x"e408902b",
  2465 => x"83fff00a",
  2466 => x"06707507",
  2467 => x"51537280",
  2468 => x"ef800c80",
  2469 => x"ef800853",
  2470 => x"72802e9e",
  2471 => x"3880eed4",
  2472 => x"08fe1471",
  2473 => x"2980eee8",
  2474 => x"080580ef",
  2475 => x"840c7084",
  2476 => x"2b80eee0",
  2477 => x"0c5480cd",
  2478 => x"e90480ee",
  2479 => x"ec0880ef",
  2480 => x"800c80ee",
  2481 => x"f00880ef",
  2482 => x"840c80ee",
  2483 => x"dc08802e",
  2484 => x"8c3880ee",
  2485 => x"d408842b",
  2486 => x"5380cde4",
  2487 => x"0480eef4",
  2488 => x"08842b53",
  2489 => x"7280eee0",
  2490 => x"0c029405",
  2491 => x"0d0402d8",
  2492 => x"050d800b",
  2493 => x"80eedc0c",
  2494 => x"845480c7",
  2495 => x"c72d80e7",
  2496 => x"e408802e",
  2497 => x"993880e8",
  2498 => x"d0528051",
  2499 => x"80cadb2d",
  2500 => x"80e7e408",
  2501 => x"802e8738",
  2502 => x"fe5480ce",
  2503 => x"a604ff14",
  2504 => x"54738024",
  2505 => x"d538738e",
  2506 => x"3880e3b0",
  2507 => x"5186a02d",
  2508 => x"735580d4",
  2509 => x"8a048056",
  2510 => x"810b80ef",
  2511 => x"880c8853",
  2512 => x"80e3c452",
  2513 => x"80e98651",
  2514 => x"80cc832d",
  2515 => x"80e7e408",
  2516 => x"762e0981",
  2517 => x"06893880",
  2518 => x"e7e40880",
  2519 => x"ef880c88",
  2520 => x"5380e3d0",
  2521 => x"5280e9a2",
  2522 => x"5180cc83",
  2523 => x"2d80e7e4",
  2524 => x"08893880",
  2525 => x"e7e40880",
  2526 => x"ef880c80",
  2527 => x"ef880880",
  2528 => x"2e818538",
  2529 => x"80ec960b",
  2530 => x"80f52d80",
  2531 => x"ec970b80",
  2532 => x"f52d7198",
  2533 => x"2b71902b",
  2534 => x"0780ec98",
  2535 => x"0b80f52d",
  2536 => x"70882b72",
  2537 => x"0780ec99",
  2538 => x"0b80f52d",
  2539 => x"710780ec",
  2540 => x"ce0b80f5",
  2541 => x"2d80eccf",
  2542 => x"0b80f52d",
  2543 => x"71882b07",
  2544 => x"535f5452",
  2545 => x"5a565755",
  2546 => x"7381abaa",
  2547 => x"2e098106",
  2548 => x"90387551",
  2549 => x"80dace2d",
  2550 => x"80e7e408",
  2551 => x"5680cff0",
  2552 => x"047382d4",
  2553 => x"d52e8938",
  2554 => x"80e3dc51",
  2555 => x"80d0c004",
  2556 => x"80e8d052",
  2557 => x"755180ca",
  2558 => x"db2d80e7",
  2559 => x"e4085580",
  2560 => x"e7e40880",
  2561 => x"2e848338",
  2562 => x"885380e3",
  2563 => x"d05280e9",
  2564 => x"a25180cc",
  2565 => x"832d80e7",
  2566 => x"e4088b38",
  2567 => x"810b80ee",
  2568 => x"dc0c80d0",
  2569 => x"c7048853",
  2570 => x"80e3c452",
  2571 => x"80e98651",
  2572 => x"80cc832d",
  2573 => x"80e7e408",
  2574 => x"802e8c38",
  2575 => x"80e3f051",
  2576 => x"86a02d80",
  2577 => x"d1a60480",
  2578 => x"ecce0b80",
  2579 => x"f52d5473",
  2580 => x"80d52e09",
  2581 => x"810680ce",
  2582 => x"3880eccf",
  2583 => x"0b80f52d",
  2584 => x"547381aa",
  2585 => x"2e098106",
  2586 => x"bd38800b",
  2587 => x"80e8d00b",
  2588 => x"80f52d56",
  2589 => x"547481e9",
  2590 => x"2e833881",
  2591 => x"547481eb",
  2592 => x"2e8c3880",
  2593 => x"5573752e",
  2594 => x"09810682",
  2595 => x"fd3880e8",
  2596 => x"db0b80f5",
  2597 => x"2d55748e",
  2598 => x"3880e8dc",
  2599 => x"0b80f52d",
  2600 => x"5473822e",
  2601 => x"87388055",
  2602 => x"80d48a04",
  2603 => x"80e8dd0b",
  2604 => x"80f52d70",
  2605 => x"80eed40c",
  2606 => x"ff0580ee",
  2607 => x"d80c80e8",
  2608 => x"de0b80f5",
  2609 => x"2d80e8df",
  2610 => x"0b80f52d",
  2611 => x"58760577",
  2612 => x"82802905",
  2613 => x"7080eee4",
  2614 => x"0c80e8e0",
  2615 => x"0b80f52d",
  2616 => x"7080eef8",
  2617 => x"0c80eedc",
  2618 => x"08595758",
  2619 => x"76802e81",
  2620 => x"b9388853",
  2621 => x"80e3d052",
  2622 => x"80e9a251",
  2623 => x"80cc832d",
  2624 => x"80e7e408",
  2625 => x"82843880",
  2626 => x"eed40870",
  2627 => x"842b80ee",
  2628 => x"e00c7080",
  2629 => x"eef40c80",
  2630 => x"e8f50b80",
  2631 => x"f52d80e8",
  2632 => x"f40b80f5",
  2633 => x"2d718280",
  2634 => x"290580e8",
  2635 => x"f60b80f5",
  2636 => x"2d708480",
  2637 => x"80291280",
  2638 => x"e8f70b80",
  2639 => x"f52d7081",
  2640 => x"800a2912",
  2641 => x"7080eefc",
  2642 => x"0c80eef8",
  2643 => x"08712980",
  2644 => x"eee40805",
  2645 => x"7080eee8",
  2646 => x"0c80e8fd",
  2647 => x"0b80f52d",
  2648 => x"80e8fc0b",
  2649 => x"80f52d71",
  2650 => x"82802905",
  2651 => x"80e8fe0b",
  2652 => x"80f52d70",
  2653 => x"84808029",
  2654 => x"1280e8ff",
  2655 => x"0b80f52d",
  2656 => x"70982b81",
  2657 => x"f00a0672",
  2658 => x"057080ee",
  2659 => x"ec0cfe11",
  2660 => x"7e297705",
  2661 => x"80eef00c",
  2662 => x"52595243",
  2663 => x"545e5152",
  2664 => x"59525d57",
  2665 => x"595780d4",
  2666 => x"820480e8",
  2667 => x"e20b80f5",
  2668 => x"2d80e8e1",
  2669 => x"0b80f52d",
  2670 => x"71828029",
  2671 => x"057080ee",
  2672 => x"e00c70a0",
  2673 => x"2983ff05",
  2674 => x"70892a70",
  2675 => x"80eef40c",
  2676 => x"80e8e70b",
  2677 => x"80f52d80",
  2678 => x"e8e60b80",
  2679 => x"f52d7182",
  2680 => x"80290570",
  2681 => x"80eefc0c",
  2682 => x"7b71291e",
  2683 => x"7080eef0",
  2684 => x"0c7d80ee",
  2685 => x"ec0c7305",
  2686 => x"80eee80c",
  2687 => x"555e5151",
  2688 => x"55558051",
  2689 => x"80ccc42d",
  2690 => x"81557480",
  2691 => x"e7e40c02",
  2692 => x"a8050d04",
  2693 => x"02ec050d",
  2694 => x"7670872c",
  2695 => x"7180ff06",
  2696 => x"55565480",
  2697 => x"eedc088a",
  2698 => x"3873882c",
  2699 => x"7481ff06",
  2700 => x"545580e8",
  2701 => x"d05280ee",
  2702 => x"e4081551",
  2703 => x"80cadb2d",
  2704 => x"80e7e408",
  2705 => x"5480e7e4",
  2706 => x"08802ebb",
  2707 => x"3880eedc",
  2708 => x"08802e9c",
  2709 => x"38728429",
  2710 => x"80e8d005",
  2711 => x"70085253",
  2712 => x"80dace2d",
  2713 => x"80e7e408",
  2714 => x"f00a0653",
  2715 => x"80d58504",
  2716 => x"721080e8",
  2717 => x"d0057080",
  2718 => x"e02d5253",
  2719 => x"80daff2d",
  2720 => x"80e7e408",
  2721 => x"53725473",
  2722 => x"80e7e40c",
  2723 => x"0294050d",
  2724 => x"0402e005",
  2725 => x"0d797084",
  2726 => x"2c80ef84",
  2727 => x"0805718f",
  2728 => x"06525553",
  2729 => x"728b3880",
  2730 => x"e8d05273",
  2731 => x"5180cadb",
  2732 => x"2d72a029",
  2733 => x"80e8d005",
  2734 => x"54807480",
  2735 => x"f52d5653",
  2736 => x"74732e83",
  2737 => x"38815374",
  2738 => x"81e52e81",
  2739 => x"f5388170",
  2740 => x"74065458",
  2741 => x"72802e81",
  2742 => x"e9388b14",
  2743 => x"80f52d70",
  2744 => x"832a7906",
  2745 => x"5856769c",
  2746 => x"3880e6a8",
  2747 => x"08537289",
  2748 => x"387280ec",
  2749 => x"d00b81b7",
  2750 => x"2d7680e6",
  2751 => x"a80c7353",
  2752 => x"80d7c404",
  2753 => x"758f2e09",
  2754 => x"810681b6",
  2755 => x"38749f06",
  2756 => x"8d2980ec",
  2757 => x"c3115153",
  2758 => x"811480f5",
  2759 => x"2d737081",
  2760 => x"055581b7",
  2761 => x"2d831480",
  2762 => x"f52d7370",
  2763 => x"81055581",
  2764 => x"b72d8514",
  2765 => x"80f52d73",
  2766 => x"70810555",
  2767 => x"81b72d87",
  2768 => x"1480f52d",
  2769 => x"73708105",
  2770 => x"5581b72d",
  2771 => x"891480f5",
  2772 => x"2d737081",
  2773 => x"055581b7",
  2774 => x"2d8e1480",
  2775 => x"f52d7370",
  2776 => x"81055581",
  2777 => x"b72d9014",
  2778 => x"80f52d73",
  2779 => x"70810555",
  2780 => x"81b72d92",
  2781 => x"1480f52d",
  2782 => x"73708105",
  2783 => x"5581b72d",
  2784 => x"941480f5",
  2785 => x"2d737081",
  2786 => x"055581b7",
  2787 => x"2d961480",
  2788 => x"f52d7370",
  2789 => x"81055581",
  2790 => x"b72d9814",
  2791 => x"80f52d73",
  2792 => x"70810555",
  2793 => x"81b72d9c",
  2794 => x"1480f52d",
  2795 => x"73708105",
  2796 => x"5581b72d",
  2797 => x"9e1480f5",
  2798 => x"2d7381b7",
  2799 => x"2d7780e6",
  2800 => x"a80c8053",
  2801 => x"7280e7e4",
  2802 => x"0c02a005",
  2803 => x"0d0402cc",
  2804 => x"050d7e60",
  2805 => x"5e5a800b",
  2806 => x"80ef8008",
  2807 => x"80ef8408",
  2808 => x"595c5680",
  2809 => x"5880eee0",
  2810 => x"08782e81",
  2811 => x"be38778f",
  2812 => x"06a01757",
  2813 => x"54739238",
  2814 => x"80e8d052",
  2815 => x"76518117",
  2816 => x"5780cadb",
  2817 => x"2d80e8d0",
  2818 => x"56807680",
  2819 => x"f52d5654",
  2820 => x"74742e83",
  2821 => x"38815474",
  2822 => x"81e52e81",
  2823 => x"82388170",
  2824 => x"7506555c",
  2825 => x"73802e80",
  2826 => x"f6388b16",
  2827 => x"80f52d98",
  2828 => x"06597880",
  2829 => x"ea388b53",
  2830 => x"7c527551",
  2831 => x"80cc832d",
  2832 => x"80e7e408",
  2833 => x"80d9389c",
  2834 => x"16085180",
  2835 => x"dace2d80",
  2836 => x"e7e40884",
  2837 => x"1b0c9a16",
  2838 => x"80e02d51",
  2839 => x"80daff2d",
  2840 => x"80e7e408",
  2841 => x"80e7e408",
  2842 => x"881c0c80",
  2843 => x"e7e40855",
  2844 => x"5580eedc",
  2845 => x"08802e9a",
  2846 => x"38941680",
  2847 => x"e02d5180",
  2848 => x"daff2d80",
  2849 => x"e7e40890",
  2850 => x"2b83fff0",
  2851 => x"0a067016",
  2852 => x"51547388",
  2853 => x"1b0c787a",
  2854 => x"0c7b5480",
  2855 => x"d9e90481",
  2856 => x"185880ee",
  2857 => x"e0087826",
  2858 => x"fec43880",
  2859 => x"eedc0880",
  2860 => x"2eb5387a",
  2861 => x"5180d494",
  2862 => x"2d80e7e4",
  2863 => x"0880e7e4",
  2864 => x"0880ffff",
  2865 => x"fff80655",
  2866 => x"5b7380ff",
  2867 => x"fffff82e",
  2868 => x"963880e7",
  2869 => x"e408fe05",
  2870 => x"80eed408",
  2871 => x"2980eee8",
  2872 => x"08055780",
  2873 => x"d7e30480",
  2874 => x"547380e7",
  2875 => x"e40c02b4",
  2876 => x"050d0402",
  2877 => x"f4050d74",
  2878 => x"70088105",
  2879 => x"710c7008",
  2880 => x"80eed808",
  2881 => x"06535371",
  2882 => x"90388813",
  2883 => x"085180d4",
  2884 => x"942d80e7",
  2885 => x"e4088814",
  2886 => x"0c810b80",
  2887 => x"e7e40c02",
  2888 => x"8c050d04",
  2889 => x"02f0050d",
  2890 => x"75881108",
  2891 => x"fe0580ee",
  2892 => x"d4082980",
  2893 => x"eee80811",
  2894 => x"720880ee",
  2895 => x"d8080605",
  2896 => x"79555354",
  2897 => x"5480cadb",
  2898 => x"2d029005",
  2899 => x"0d0402f4",
  2900 => x"050d7470",
  2901 => x"882a83fe",
  2902 => x"80067072",
  2903 => x"982a0772",
  2904 => x"882b87fc",
  2905 => x"80800673",
  2906 => x"982b81f0",
  2907 => x"0a067173",
  2908 => x"070780e7",
  2909 => x"e40c5651",
  2910 => x"5351028c",
  2911 => x"050d0402",
  2912 => x"f8050d02",
  2913 => x"8e0580f5",
  2914 => x"2d74882b",
  2915 => x"077083ff",
  2916 => x"ff0680e7",
  2917 => x"e40c5102",
  2918 => x"88050d04",
  2919 => x"02f4050d",
  2920 => x"74767853",
  2921 => x"54528071",
  2922 => x"25973872",
  2923 => x"70810554",
  2924 => x"80f52d72",
  2925 => x"70810554",
  2926 => x"81b72dff",
  2927 => x"115170eb",
  2928 => x"38807281",
  2929 => x"b72d028c",
  2930 => x"050d0402",
  2931 => x"e8050d77",
  2932 => x"56807056",
  2933 => x"54737624",
  2934 => x"b73880ee",
  2935 => x"e008742e",
  2936 => x"af387351",
  2937 => x"80d5912d",
  2938 => x"80e7e408",
  2939 => x"80e7e408",
  2940 => x"09810570",
  2941 => x"80e7e408",
  2942 => x"079f2a77",
  2943 => x"05811757",
  2944 => x"57535374",
  2945 => x"76248938",
  2946 => x"80eee008",
  2947 => x"7426d338",
  2948 => x"7280e7e4",
  2949 => x"0c029805",
  2950 => x"0d0402f0",
  2951 => x"050d80e7",
  2952 => x"e0081651",
  2953 => x"80dbcb2d",
  2954 => x"80e7e408",
  2955 => x"802ea038",
  2956 => x"8b5380e7",
  2957 => x"e4085280",
  2958 => x"ecd05180",
  2959 => x"db9c2d80",
  2960 => x"ef8c0854",
  2961 => x"73802e87",
  2962 => x"3880ecd0",
  2963 => x"51732d02",
  2964 => x"90050d04",
  2965 => x"02dc050d",
  2966 => x"80705a55",
  2967 => x"7480e7e0",
  2968 => x"0825b538",
  2969 => x"80eee008",
  2970 => x"752ead38",
  2971 => x"785180d5",
  2972 => x"912d80e7",
  2973 => x"e4080981",
  2974 => x"057080e7",
  2975 => x"e408079f",
  2976 => x"2a760581",
  2977 => x"1b5b5654",
  2978 => x"7480e7e0",
  2979 => x"08258938",
  2980 => x"80eee008",
  2981 => x"7926d538",
  2982 => x"80557880",
  2983 => x"eee00827",
  2984 => x"81e43878",
  2985 => x"5180d591",
  2986 => x"2d80e7e4",
  2987 => x"08802e81",
  2988 => x"b43880e7",
  2989 => x"e4088b05",
  2990 => x"80f52d70",
  2991 => x"842a7081",
  2992 => x"06771078",
  2993 => x"842b80ec",
  2994 => x"d00b80f5",
  2995 => x"2d5c5c53",
  2996 => x"51555673",
  2997 => x"802e80ce",
  2998 => x"38741682",
  2999 => x"2b80dfaa",
  3000 => x"0b80e6b4",
  3001 => x"120c5477",
  3002 => x"75311080",
  3003 => x"ef901155",
  3004 => x"56907470",
  3005 => x"81055681",
  3006 => x"b72da074",
  3007 => x"81b72d76",
  3008 => x"81ff0681",
  3009 => x"16585473",
  3010 => x"802e8b38",
  3011 => x"9c5380ec",
  3012 => x"d05280de",
  3013 => x"9d048b53",
  3014 => x"80e7e408",
  3015 => x"5280ef92",
  3016 => x"165180de",
  3017 => x"db047416",
  3018 => x"822b80dc",
  3019 => x"9a0b80e6",
  3020 => x"b4120c54",
  3021 => x"7681ff06",
  3022 => x"81165854",
  3023 => x"73802e8b",
  3024 => x"389c5380",
  3025 => x"ecd05280",
  3026 => x"ded2048b",
  3027 => x"5380e7e4",
  3028 => x"08527775",
  3029 => x"311080ef",
  3030 => x"90055176",
  3031 => x"5580db9c",
  3032 => x"2d80defa",
  3033 => x"04749029",
  3034 => x"75317010",
  3035 => x"80ef9005",
  3036 => x"515480e7",
  3037 => x"e4087481",
  3038 => x"b72d8119",
  3039 => x"59748b24",
  3040 => x"a43880dd",
  3041 => x"9a047490",
  3042 => x"29753170",
  3043 => x"1080ef90",
  3044 => x"058c7731",
  3045 => x"57515480",
  3046 => x"7481b72d",
  3047 => x"9e14ff16",
  3048 => x"565474f3",
  3049 => x"3802a405",
  3050 => x"0d0402fc",
  3051 => x"050d80e7",
  3052 => x"e0081351",
  3053 => x"80dbcb2d",
  3054 => x"80e7e408",
  3055 => x"802e8a38",
  3056 => x"80e7e408",
  3057 => x"5180ccc4",
  3058 => x"2d800b80",
  3059 => x"e7e00c80",
  3060 => x"dcd42db9",
  3061 => x"d42d0284",
  3062 => x"050d0402",
  3063 => x"fc050d72",
  3064 => x"5170fd2e",
  3065 => x"b23870fd",
  3066 => x"248b3870",
  3067 => x"fc2e80d0",
  3068 => x"3880e0ca",
  3069 => x"0470fe2e",
  3070 => x"b93870ff",
  3071 => x"2e098106",
  3072 => x"80c83880",
  3073 => x"e7e00851",
  3074 => x"70802ebe",
  3075 => x"38ff1180",
  3076 => x"e7e00c80",
  3077 => x"e0ca0480",
  3078 => x"e7e008f0",
  3079 => x"057080e7",
  3080 => x"e00c5170",
  3081 => x"8025a338",
  3082 => x"800b80e7",
  3083 => x"e00c80e0",
  3084 => x"ca0480e7",
  3085 => x"e0088105",
  3086 => x"80e7e00c",
  3087 => x"80e0ca04",
  3088 => x"80e7e008",
  3089 => x"900580e7",
  3090 => x"e00c80dc",
  3091 => x"d42db9d4",
  3092 => x"2d028405",
  3093 => x"0d0402fc",
  3094 => x"050d800b",
  3095 => x"80e7e00c",
  3096 => x"80dcd42d",
  3097 => x"b8c22d80",
  3098 => x"e7e40880",
  3099 => x"e7d00c80",
  3100 => x"e6ac51ba",
  3101 => x"fa2d0284",
  3102 => x"050d0471",
  3103 => x"80ef8c0c",
  3104 => x"04000000",
  3105 => x"00ffffff",
  3106 => x"ff00ffff",
  3107 => x"ffff00ff",
  3108 => x"ffffff00",
  3109 => x"4b455953",
  3110 => x"50312020",
  3111 => x"20202000",
  3112 => x"00000000",
  3113 => x"4b455953",
  3114 => x"50322020",
  3115 => x"20202000",
  3116 => x"00000000",
  3117 => x"52657365",
  3118 => x"74000000",
  3119 => x"5363616e",
  3120 => x"6c696e65",
  3121 => x"73000000",
  3122 => x"50414c20",
  3123 => x"2f204e54",
  3124 => x"53430000",
  3125 => x"436f6c6f",
  3126 => x"72000000",
  3127 => x"44696666",
  3128 => x"6963756c",
  3129 => x"74792041",
  3130 => x"00000000",
  3131 => x"44696666",
  3132 => x"6963756c",
  3133 => x"74792042",
  3134 => x"00000000",
  3135 => x"53656c65",
  3136 => x"63740000",
  3137 => x"53746172",
  3138 => x"74000000",
  3139 => x"4c6f6164",
  3140 => x"20524f4d",
  3141 => x"20100000",
  3142 => x"45786974",
  3143 => x"00000000",
  3144 => x"524f4d20",
  3145 => x"6c6f6164",
  3146 => x"696e6720",
  3147 => x"6661696c",
  3148 => x"65640000",
  3149 => x"4f4b0000",
  3150 => x"496e6974",
  3151 => x"69616c69",
  3152 => x"7a696e67",
  3153 => x"20534420",
  3154 => x"63617264",
  3155 => x"0a000000",
  3156 => x"16200000",
  3157 => x"14200000",
  3158 => x"15200000",
  3159 => x"53442069",
  3160 => x"6e69742e",
  3161 => x"2e2e0a00",
  3162 => x"53442063",
  3163 => x"61726420",
  3164 => x"72657365",
  3165 => x"74206661",
  3166 => x"696c6564",
  3167 => x"210a0000",
  3168 => x"53444843",
  3169 => x"20657272",
  3170 => x"6f72210a",
  3171 => x"00000000",
  3172 => x"57726974",
  3173 => x"65206661",
  3174 => x"696c6564",
  3175 => x"0a000000",
  3176 => x"52656164",
  3177 => x"20666169",
  3178 => x"6c65640a",
  3179 => x"00000000",
  3180 => x"43617264",
  3181 => x"20696e69",
  3182 => x"74206661",
  3183 => x"696c6564",
  3184 => x"0a000000",
  3185 => x"46415431",
  3186 => x"36202020",
  3187 => x"00000000",
  3188 => x"46415433",
  3189 => x"32202020",
  3190 => x"00000000",
  3191 => x"4e6f2070",
  3192 => x"61727469",
  3193 => x"74696f6e",
  3194 => x"20736967",
  3195 => x"0a000000",
  3196 => x"42616420",
  3197 => x"70617274",
  3198 => x"0a000000",
  3199 => x"4261636b",
  3200 => x"00000000",
  3201 => x"00000002",
  3202 => x"00000002",
  3203 => x"000030b4",
  3204 => x"0000035a",
  3205 => x"00000001",
  3206 => x"000030bc",
  3207 => x"00000000",
  3208 => x"00000001",
  3209 => x"000030c8",
  3210 => x"00000001",
  3211 => x"00000001",
  3212 => x"000030d4",
  3213 => x"00000002",
  3214 => x"00000001",
  3215 => x"000030dc",
  3216 => x"00000003",
  3217 => x"00000001",
  3218 => x"000030ec",
  3219 => x"00000004",
  3220 => x"00000002",
  3221 => x"000030fc",
  3222 => x"0000036e",
  3223 => x"00000002",
  3224 => x"00003104",
  3225 => x"00000a3f",
  3226 => x"00000002",
  3227 => x"0000310c",
  3228 => x"00003056",
  3229 => x"00000002",
  3230 => x"00003118",
  3231 => x"00001c5f",
  3232 => x"00000000",
  3233 => x"00000000",
  3234 => x"00000000",
  3235 => x"00000004",
  3236 => x"00003120",
  3237 => x"0000328c",
  3238 => x"00000004",
  3239 => x"00003134",
  3240 => x"00003208",
  3241 => x"00000000",
  3242 => x"00000000",
  3243 => x"00000000",
  3244 => x"00000000",
  3245 => x"00000000",
  3246 => x"00000000",
  3247 => x"00000000",
  3248 => x"00000000",
  3249 => x"00000000",
  3250 => x"00000000",
  3251 => x"00000000",
  3252 => x"00000000",
  3253 => x"00000000",
  3254 => x"00000000",
  3255 => x"00000000",
  3256 => x"00000000",
  3257 => x"00000000",
  3258 => x"00000000",
  3259 => x"00000000",
  3260 => x"00000000",
  3261 => x"00000000",
  3262 => x"00000006",
  3263 => x"00000043",
  3264 => x"00000042",
  3265 => x"0000003b",
  3266 => x"0000004b",
  3267 => x"00000033",
  3268 => x"0000001d",
  3269 => x"0000001b",
  3270 => x"0000001c",
  3271 => x"00000023",
  3272 => x"0000002b",
  3273 => x"00000000",
  3274 => x"00000000",
  3275 => x"00000002",
  3276 => x"00003790",
  3277 => x"00002e1a",
  3278 => x"00000002",
  3279 => x"000037ae",
  3280 => x"00002e1a",
  3281 => x"00000002",
  3282 => x"000037cc",
  3283 => x"00002e1a",
  3284 => x"00000002",
  3285 => x"000037ea",
  3286 => x"00002e1a",
  3287 => x"00000002",
  3288 => x"00003808",
  3289 => x"00002e1a",
  3290 => x"00000002",
  3291 => x"00003826",
  3292 => x"00002e1a",
  3293 => x"00000002",
  3294 => x"00003844",
  3295 => x"00002e1a",
  3296 => x"00000002",
  3297 => x"00003862",
  3298 => x"00002e1a",
  3299 => x"00000002",
  3300 => x"00003880",
  3301 => x"00002e1a",
  3302 => x"00000002",
  3303 => x"0000389e",
  3304 => x"00002e1a",
  3305 => x"00000002",
  3306 => x"000038bc",
  3307 => x"00002e1a",
  3308 => x"00000002",
  3309 => x"000038da",
  3310 => x"00002e1a",
  3311 => x"00000002",
  3312 => x"000038f8",
  3313 => x"00002e1a",
  3314 => x"00000004",
  3315 => x"000031fc",
  3316 => x"00000000",
  3317 => x"00000000",
  3318 => x"00000000",
  3319 => x"00002fdb",
  3320 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

